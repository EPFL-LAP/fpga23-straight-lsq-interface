module STORE_QUEUE_LSQ_data( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input         io_bbStart, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_0, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_1, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_2, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_3, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_4, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_5, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_6, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_7, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_8, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_9, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_10, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_11, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_12, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_13, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_14, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_15, // @[:@6.4]
  input  [1:0]  io_bbNumStores, // @[:@6.4]
  output [3:0]  io_storeTail, // @[:@6.4]
  output [3:0]  io_storeHead, // @[:@6.4]
  output        io_storeEmpty, // @[:@6.4]
  input  [3:0]  io_loadTail, // @[:@6.4]
  input  [3:0]  io_loadHead, // @[:@6.4]
  input         io_loadEmpty, // @[:@6.4]
  input         io_loadAddressDone_0, // @[:@6.4]
  input         io_loadAddressDone_1, // @[:@6.4]
  input         io_loadAddressDone_2, // @[:@6.4]
  input         io_loadAddressDone_3, // @[:@6.4]
  input         io_loadAddressDone_4, // @[:@6.4]
  input         io_loadAddressDone_5, // @[:@6.4]
  input         io_loadAddressDone_6, // @[:@6.4]
  input         io_loadAddressDone_7, // @[:@6.4]
  input         io_loadAddressDone_8, // @[:@6.4]
  input         io_loadAddressDone_9, // @[:@6.4]
  input         io_loadAddressDone_10, // @[:@6.4]
  input         io_loadAddressDone_11, // @[:@6.4]
  input         io_loadAddressDone_12, // @[:@6.4]
  input         io_loadAddressDone_13, // @[:@6.4]
  input         io_loadAddressDone_14, // @[:@6.4]
  input         io_loadAddressDone_15, // @[:@6.4]
  input         io_loadDataDone_0, // @[:@6.4]
  input         io_loadDataDone_1, // @[:@6.4]
  input         io_loadDataDone_2, // @[:@6.4]
  input         io_loadDataDone_3, // @[:@6.4]
  input         io_loadDataDone_4, // @[:@6.4]
  input         io_loadDataDone_5, // @[:@6.4]
  input         io_loadDataDone_6, // @[:@6.4]
  input         io_loadDataDone_7, // @[:@6.4]
  input         io_loadDataDone_8, // @[:@6.4]
  input         io_loadDataDone_9, // @[:@6.4]
  input         io_loadDataDone_10, // @[:@6.4]
  input         io_loadDataDone_11, // @[:@6.4]
  input         io_loadDataDone_12, // @[:@6.4]
  input         io_loadDataDone_13, // @[:@6.4]
  input         io_loadDataDone_14, // @[:@6.4]
  input         io_loadDataDone_15, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_0, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_1, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_2, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_3, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_4, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_5, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_6, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_7, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_8, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_9, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_10, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_11, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_12, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_13, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_14, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_15, // @[:@6.4]
  output        io_storeAddrDone_0, // @[:@6.4]
  output        io_storeAddrDone_1, // @[:@6.4]
  output        io_storeAddrDone_2, // @[:@6.4]
  output        io_storeAddrDone_3, // @[:@6.4]
  output        io_storeAddrDone_4, // @[:@6.4]
  output        io_storeAddrDone_5, // @[:@6.4]
  output        io_storeAddrDone_6, // @[:@6.4]
  output        io_storeAddrDone_7, // @[:@6.4]
  output        io_storeAddrDone_8, // @[:@6.4]
  output        io_storeAddrDone_9, // @[:@6.4]
  output        io_storeAddrDone_10, // @[:@6.4]
  output        io_storeAddrDone_11, // @[:@6.4]
  output        io_storeAddrDone_12, // @[:@6.4]
  output        io_storeAddrDone_13, // @[:@6.4]
  output        io_storeAddrDone_14, // @[:@6.4]
  output        io_storeAddrDone_15, // @[:@6.4]
  output        io_storeDataDone_0, // @[:@6.4]
  output        io_storeDataDone_1, // @[:@6.4]
  output        io_storeDataDone_2, // @[:@6.4]
  output        io_storeDataDone_3, // @[:@6.4]
  output        io_storeDataDone_4, // @[:@6.4]
  output        io_storeDataDone_5, // @[:@6.4]
  output        io_storeDataDone_6, // @[:@6.4]
  output        io_storeDataDone_7, // @[:@6.4]
  output        io_storeDataDone_8, // @[:@6.4]
  output        io_storeDataDone_9, // @[:@6.4]
  output        io_storeDataDone_10, // @[:@6.4]
  output        io_storeDataDone_11, // @[:@6.4]
  output        io_storeDataDone_12, // @[:@6.4]
  output        io_storeDataDone_13, // @[:@6.4]
  output        io_storeDataDone_14, // @[:@6.4]
  output        io_storeDataDone_15, // @[:@6.4]
  output [31:0] io_storeAddrQueue_0, // @[:@6.4]
  output [31:0] io_storeAddrQueue_1, // @[:@6.4]
  output [31:0] io_storeAddrQueue_2, // @[:@6.4]
  output [31:0] io_storeAddrQueue_3, // @[:@6.4]
  output [31:0] io_storeAddrQueue_4, // @[:@6.4]
  output [31:0] io_storeAddrQueue_5, // @[:@6.4]
  output [31:0] io_storeAddrQueue_6, // @[:@6.4]
  output [31:0] io_storeAddrQueue_7, // @[:@6.4]
  output [31:0] io_storeAddrQueue_8, // @[:@6.4]
  output [31:0] io_storeAddrQueue_9, // @[:@6.4]
  output [31:0] io_storeAddrQueue_10, // @[:@6.4]
  output [31:0] io_storeAddrQueue_11, // @[:@6.4]
  output [31:0] io_storeAddrQueue_12, // @[:@6.4]
  output [31:0] io_storeAddrQueue_13, // @[:@6.4]
  output [31:0] io_storeAddrQueue_14, // @[:@6.4]
  output [31:0] io_storeAddrQueue_15, // @[:@6.4]
  output [31:0] io_storeDataQueue_0, // @[:@6.4]
  output [31:0] io_storeDataQueue_1, // @[:@6.4]
  output [31:0] io_storeDataQueue_2, // @[:@6.4]
  output [31:0] io_storeDataQueue_3, // @[:@6.4]
  output [31:0] io_storeDataQueue_4, // @[:@6.4]
  output [31:0] io_storeDataQueue_5, // @[:@6.4]
  output [31:0] io_storeDataQueue_6, // @[:@6.4]
  output [31:0] io_storeDataQueue_7, // @[:@6.4]
  output [31:0] io_storeDataQueue_8, // @[:@6.4]
  output [31:0] io_storeDataQueue_9, // @[:@6.4]
  output [31:0] io_storeDataQueue_10, // @[:@6.4]
  output [31:0] io_storeDataQueue_11, // @[:@6.4]
  output [31:0] io_storeDataQueue_12, // @[:@6.4]
  output [31:0] io_storeDataQueue_13, // @[:@6.4]
  output [31:0] io_storeDataQueue_14, // @[:@6.4]
  output [31:0] io_storeDataQueue_15, // @[:@6.4]
  input         io_storeDataEnable_0, // @[:@6.4]
  input  [31:0] io_dataFromStorePorts_0, // @[:@6.4]
  input         io_storeAddrEnable_0, // @[:@6.4]
  input  [31:0] io_addressFromStorePorts_0, // @[:@6.4]
  output [31:0] io_storeAddrToMem, // @[:@6.4]
  output [31:0] io_storeDataToMem, // @[:@6.4]
  output        io_storeEnableToMem, // @[:@6.4]
  input         io_memIsReadyForStores // @[:@6.4]
);
  reg [3:0] head; // @[StoreQueue.scala 50:21:@8.4]
  reg [31:0] _RAND_0;
  reg [3:0] tail; // @[StoreQueue.scala 51:21:@9.4]
  reg [31:0] _RAND_1;
  reg [3:0] offsetQ_0; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_2;
  reg [3:0] offsetQ_1; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_3;
  reg [3:0] offsetQ_2; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_4;
  reg [3:0] offsetQ_3; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_5;
  reg [3:0] offsetQ_4; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_6;
  reg [3:0] offsetQ_5; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_7;
  reg [3:0] offsetQ_6; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_8;
  reg [3:0] offsetQ_7; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_9;
  reg [3:0] offsetQ_8; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_10;
  reg [3:0] offsetQ_9; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_11;
  reg [3:0] offsetQ_10; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_12;
  reg [3:0] offsetQ_11; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_13;
  reg [3:0] offsetQ_12; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_14;
  reg [3:0] offsetQ_13; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_15;
  reg [3:0] offsetQ_14; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_16;
  reg [3:0] offsetQ_15; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_17;
  reg  portQ_0; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_18;
  reg  portQ_1; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_19;
  reg  portQ_2; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_20;
  reg  portQ_3; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_21;
  reg  portQ_4; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_22;
  reg  portQ_5; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_23;
  reg  portQ_6; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_24;
  reg  portQ_7; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_25;
  reg  portQ_8; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_26;
  reg  portQ_9; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_27;
  reg  portQ_10; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_28;
  reg  portQ_11; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_29;
  reg  portQ_12; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_30;
  reg  portQ_13; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_31;
  reg  portQ_14; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_32;
  reg  portQ_15; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_33;
  reg [31:0] addrQ_0; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_34;
  reg [31:0] addrQ_1; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_35;
  reg [31:0] addrQ_2; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_36;
  reg [31:0] addrQ_3; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_37;
  reg [31:0] addrQ_4; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_38;
  reg [31:0] addrQ_5; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_39;
  reg [31:0] addrQ_6; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_40;
  reg [31:0] addrQ_7; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_41;
  reg [31:0] addrQ_8; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_42;
  reg [31:0] addrQ_9; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_43;
  reg [31:0] addrQ_10; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_44;
  reg [31:0] addrQ_11; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_45;
  reg [31:0] addrQ_12; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_46;
  reg [31:0] addrQ_13; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_47;
  reg [31:0] addrQ_14; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_48;
  reg [31:0] addrQ_15; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_49;
  reg [31:0] dataQ_0; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_50;
  reg [31:0] dataQ_1; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_51;
  reg [31:0] dataQ_2; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_52;
  reg [31:0] dataQ_3; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_53;
  reg [31:0] dataQ_4; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_54;
  reg [31:0] dataQ_5; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_55;
  reg [31:0] dataQ_6; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_56;
  reg [31:0] dataQ_7; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_57;
  reg [31:0] dataQ_8; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_58;
  reg [31:0] dataQ_9; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_59;
  reg [31:0] dataQ_10; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_60;
  reg [31:0] dataQ_11; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_61;
  reg [31:0] dataQ_12; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_62;
  reg [31:0] dataQ_13; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_63;
  reg [31:0] dataQ_14; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_64;
  reg [31:0] dataQ_15; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_65;
  reg  addrKnown_0; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_66;
  reg  addrKnown_1; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_67;
  reg  addrKnown_2; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_68;
  reg  addrKnown_3; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_69;
  reg  addrKnown_4; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_70;
  reg  addrKnown_5; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_71;
  reg  addrKnown_6; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_72;
  reg  addrKnown_7; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_73;
  reg  addrKnown_8; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_74;
  reg  addrKnown_9; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_75;
  reg  addrKnown_10; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_76;
  reg  addrKnown_11; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_77;
  reg  addrKnown_12; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_78;
  reg  addrKnown_13; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_79;
  reg  addrKnown_14; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_80;
  reg  addrKnown_15; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_81;
  reg  dataKnown_0; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_82;
  reg  dataKnown_1; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_83;
  reg  dataKnown_2; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_84;
  reg  dataKnown_3; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_85;
  reg  dataKnown_4; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_86;
  reg  dataKnown_5; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_87;
  reg  dataKnown_6; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_88;
  reg  dataKnown_7; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_89;
  reg  dataKnown_8; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_90;
  reg  dataKnown_9; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_91;
  reg  dataKnown_10; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_92;
  reg  dataKnown_11; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_93;
  reg  dataKnown_12; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_94;
  reg  dataKnown_13; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_95;
  reg  dataKnown_14; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_96;
  reg  dataKnown_15; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_97;
  reg  allocatedEntries_0; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_98;
  reg  allocatedEntries_1; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_99;
  reg  allocatedEntries_2; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_100;
  reg  allocatedEntries_3; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_101;
  reg  allocatedEntries_4; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_102;
  reg  allocatedEntries_5; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_103;
  reg  allocatedEntries_6; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_104;
  reg  allocatedEntries_7; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_105;
  reg  allocatedEntries_8; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_106;
  reg  allocatedEntries_9; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_107;
  reg  allocatedEntries_10; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_108;
  reg  allocatedEntries_11; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_109;
  reg  allocatedEntries_12; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_110;
  reg  allocatedEntries_13; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_111;
  reg  allocatedEntries_14; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_112;
  reg  allocatedEntries_15; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_113;
  reg  storeCompleted_0; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_114;
  reg  storeCompleted_1; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_115;
  reg  storeCompleted_2; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_116;
  reg  storeCompleted_3; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_117;
  reg  storeCompleted_4; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_118;
  reg  storeCompleted_5; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_119;
  reg  storeCompleted_6; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_120;
  reg  storeCompleted_7; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_121;
  reg  storeCompleted_8; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_122;
  reg  storeCompleted_9; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_123;
  reg  storeCompleted_10; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_124;
  reg  storeCompleted_11; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_125;
  reg  storeCompleted_12; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_126;
  reg  storeCompleted_13; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_127;
  reg  storeCompleted_14; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_128;
  reg  storeCompleted_15; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_129;
  reg  checkBits_0; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_130;
  reg  checkBits_1; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_131;
  reg  checkBits_2; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_132;
  reg  checkBits_3; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_133;
  reg  checkBits_4; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_134;
  reg  checkBits_5; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_135;
  reg  checkBits_6; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_136;
  reg  checkBits_7; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_137;
  reg  checkBits_8; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_138;
  reg  checkBits_9; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_139;
  reg  checkBits_10; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_140;
  reg  checkBits_11; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_141;
  reg  checkBits_12; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_142;
  reg  checkBits_13; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_143;
  reg  checkBits_14; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_144;
  reg  checkBits_15; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_145;
  wire [5:0] _GEN_1138; // @[util.scala 14:20:@173.4]
  wire [6:0] _T_1596; // @[util.scala 14:20:@173.4]
  wire [6:0] _T_1597; // @[util.scala 14:20:@174.4]
  wire [5:0] _T_1598; // @[util.scala 14:20:@175.4]
  wire [5:0] _GEN_0; // @[util.scala 14:25:@176.4]
  wire [4:0] _T_1599; // @[util.scala 14:25:@176.4]
  wire [4:0] _GEN_1139; // @[StoreQueue.scala 70:46:@177.4]
  wire  _T_1600; // @[StoreQueue.scala 70:46:@177.4]
  wire  initBits_0; // @[StoreQueue.scala 70:64:@178.4]
  wire [6:0] _T_1605; // @[util.scala 14:20:@180.4]
  wire [6:0] _T_1606; // @[util.scala 14:20:@181.4]
  wire [5:0] _T_1607; // @[util.scala 14:20:@182.4]
  wire [5:0] _GEN_16; // @[util.scala 14:25:@183.4]
  wire [4:0] _T_1608; // @[util.scala 14:25:@183.4]
  wire  _T_1609; // @[StoreQueue.scala 70:46:@184.4]
  wire  initBits_1; // @[StoreQueue.scala 70:64:@185.4]
  wire [6:0] _T_1614; // @[util.scala 14:20:@187.4]
  wire [6:0] _T_1615; // @[util.scala 14:20:@188.4]
  wire [5:0] _T_1616; // @[util.scala 14:20:@189.4]
  wire [5:0] _GEN_17; // @[util.scala 14:25:@190.4]
  wire [4:0] _T_1617; // @[util.scala 14:25:@190.4]
  wire  _T_1618; // @[StoreQueue.scala 70:46:@191.4]
  wire  initBits_2; // @[StoreQueue.scala 70:64:@192.4]
  wire [6:0] _T_1623; // @[util.scala 14:20:@194.4]
  wire [6:0] _T_1624; // @[util.scala 14:20:@195.4]
  wire [5:0] _T_1625; // @[util.scala 14:20:@196.4]
  wire [5:0] _GEN_18; // @[util.scala 14:25:@197.4]
  wire [4:0] _T_1626; // @[util.scala 14:25:@197.4]
  wire  _T_1627; // @[StoreQueue.scala 70:46:@198.4]
  wire  initBits_3; // @[StoreQueue.scala 70:64:@199.4]
  wire [6:0] _T_1632; // @[util.scala 14:20:@201.4]
  wire [6:0] _T_1633; // @[util.scala 14:20:@202.4]
  wire [5:0] _T_1634; // @[util.scala 14:20:@203.4]
  wire [5:0] _GEN_19; // @[util.scala 14:25:@204.4]
  wire [4:0] _T_1635; // @[util.scala 14:25:@204.4]
  wire  _T_1636; // @[StoreQueue.scala 70:46:@205.4]
  wire  initBits_4; // @[StoreQueue.scala 70:64:@206.4]
  wire [6:0] _T_1641; // @[util.scala 14:20:@208.4]
  wire [6:0] _T_1642; // @[util.scala 14:20:@209.4]
  wire [5:0] _T_1643; // @[util.scala 14:20:@210.4]
  wire [5:0] _GEN_20; // @[util.scala 14:25:@211.4]
  wire [4:0] _T_1644; // @[util.scala 14:25:@211.4]
  wire  _T_1645; // @[StoreQueue.scala 70:46:@212.4]
  wire  initBits_5; // @[StoreQueue.scala 70:64:@213.4]
  wire [6:0] _T_1650; // @[util.scala 14:20:@215.4]
  wire [6:0] _T_1651; // @[util.scala 14:20:@216.4]
  wire [5:0] _T_1652; // @[util.scala 14:20:@217.4]
  wire [5:0] _GEN_21; // @[util.scala 14:25:@218.4]
  wire [4:0] _T_1653; // @[util.scala 14:25:@218.4]
  wire  _T_1654; // @[StoreQueue.scala 70:46:@219.4]
  wire  initBits_6; // @[StoreQueue.scala 70:64:@220.4]
  wire [6:0] _T_1659; // @[util.scala 14:20:@222.4]
  wire [6:0] _T_1660; // @[util.scala 14:20:@223.4]
  wire [5:0] _T_1661; // @[util.scala 14:20:@224.4]
  wire [5:0] _GEN_22; // @[util.scala 14:25:@225.4]
  wire [4:0] _T_1662; // @[util.scala 14:25:@225.4]
  wire  _T_1663; // @[StoreQueue.scala 70:46:@226.4]
  wire  initBits_7; // @[StoreQueue.scala 70:64:@227.4]
  wire [6:0] _T_1668; // @[util.scala 14:20:@229.4]
  wire [6:0] _T_1669; // @[util.scala 14:20:@230.4]
  wire [5:0] _T_1670; // @[util.scala 14:20:@231.4]
  wire [5:0] _GEN_23; // @[util.scala 14:25:@232.4]
  wire [4:0] _T_1671; // @[util.scala 14:25:@232.4]
  wire  _T_1672; // @[StoreQueue.scala 70:46:@233.4]
  wire  initBits_8; // @[StoreQueue.scala 70:64:@234.4]
  wire [6:0] _T_1677; // @[util.scala 14:20:@236.4]
  wire [6:0] _T_1678; // @[util.scala 14:20:@237.4]
  wire [5:0] _T_1679; // @[util.scala 14:20:@238.4]
  wire [5:0] _GEN_24; // @[util.scala 14:25:@239.4]
  wire [4:0] _T_1680; // @[util.scala 14:25:@239.4]
  wire  _T_1681; // @[StoreQueue.scala 70:46:@240.4]
  wire  initBits_9; // @[StoreQueue.scala 70:64:@241.4]
  wire [6:0] _T_1686; // @[util.scala 14:20:@243.4]
  wire [6:0] _T_1687; // @[util.scala 14:20:@244.4]
  wire [5:0] _T_1688; // @[util.scala 14:20:@245.4]
  wire [5:0] _GEN_25; // @[util.scala 14:25:@246.4]
  wire [4:0] _T_1689; // @[util.scala 14:25:@246.4]
  wire  _T_1690; // @[StoreQueue.scala 70:46:@247.4]
  wire  initBits_10; // @[StoreQueue.scala 70:64:@248.4]
  wire [6:0] _T_1695; // @[util.scala 14:20:@250.4]
  wire [6:0] _T_1696; // @[util.scala 14:20:@251.4]
  wire [5:0] _T_1697; // @[util.scala 14:20:@252.4]
  wire [5:0] _GEN_26; // @[util.scala 14:25:@253.4]
  wire [4:0] _T_1698; // @[util.scala 14:25:@253.4]
  wire  _T_1699; // @[StoreQueue.scala 70:46:@254.4]
  wire  initBits_11; // @[StoreQueue.scala 70:64:@255.4]
  wire [6:0] _T_1704; // @[util.scala 14:20:@257.4]
  wire [6:0] _T_1705; // @[util.scala 14:20:@258.4]
  wire [5:0] _T_1706; // @[util.scala 14:20:@259.4]
  wire [5:0] _GEN_27; // @[util.scala 14:25:@260.4]
  wire [4:0] _T_1707; // @[util.scala 14:25:@260.4]
  wire  _T_1708; // @[StoreQueue.scala 70:46:@261.4]
  wire  initBits_12; // @[StoreQueue.scala 70:64:@262.4]
  wire [6:0] _T_1713; // @[util.scala 14:20:@264.4]
  wire [6:0] _T_1714; // @[util.scala 14:20:@265.4]
  wire [5:0] _T_1715; // @[util.scala 14:20:@266.4]
  wire [5:0] _GEN_28; // @[util.scala 14:25:@267.4]
  wire [4:0] _T_1716; // @[util.scala 14:25:@267.4]
  wire  _T_1717; // @[StoreQueue.scala 70:46:@268.4]
  wire  initBits_13; // @[StoreQueue.scala 70:64:@269.4]
  wire [6:0] _T_1722; // @[util.scala 14:20:@271.4]
  wire [6:0] _T_1723; // @[util.scala 14:20:@272.4]
  wire [5:0] _T_1724; // @[util.scala 14:20:@273.4]
  wire [5:0] _GEN_29; // @[util.scala 14:25:@274.4]
  wire [4:0] _T_1725; // @[util.scala 14:25:@274.4]
  wire  _T_1726; // @[StoreQueue.scala 70:46:@275.4]
  wire  initBits_14; // @[StoreQueue.scala 70:64:@276.4]
  wire [6:0] _T_1731; // @[util.scala 14:20:@278.4]
  wire [6:0] _T_1732; // @[util.scala 14:20:@279.4]
  wire [5:0] _T_1733; // @[util.scala 14:20:@280.4]
  wire [5:0] _GEN_30; // @[util.scala 14:25:@281.4]
  wire [4:0] _T_1734; // @[util.scala 14:25:@281.4]
  wire  _T_1735; // @[StoreQueue.scala 70:46:@282.4]
  wire  initBits_15; // @[StoreQueue.scala 70:64:@283.4]
  wire  _T_1758; // @[StoreQueue.scala 72:78:@301.4]
  wire  _T_1759; // @[StoreQueue.scala 72:78:@302.4]
  wire  _T_1760; // @[StoreQueue.scala 72:78:@303.4]
  wire  _T_1761; // @[StoreQueue.scala 72:78:@304.4]
  wire  _T_1762; // @[StoreQueue.scala 72:78:@305.4]
  wire  _T_1763; // @[StoreQueue.scala 72:78:@306.4]
  wire  _T_1764; // @[StoreQueue.scala 72:78:@307.4]
  wire  _T_1765; // @[StoreQueue.scala 72:78:@308.4]
  wire  _T_1766; // @[StoreQueue.scala 72:78:@309.4]
  wire  _T_1767; // @[StoreQueue.scala 72:78:@310.4]
  wire  _T_1768; // @[StoreQueue.scala 72:78:@311.4]
  wire  _T_1769; // @[StoreQueue.scala 72:78:@312.4]
  wire  _T_1770; // @[StoreQueue.scala 72:78:@313.4]
  wire  _T_1771; // @[StoreQueue.scala 72:78:@314.4]
  wire  _T_1772; // @[StoreQueue.scala 72:78:@315.4]
  wire  _T_1773; // @[StoreQueue.scala 72:78:@316.4]
  wire [3:0] _T_1804; // @[:@356.6]
  wire [3:0] _GEN_1; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_2; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_3; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_4; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_5; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_6; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_7; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_8; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_9; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_10; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_11; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_12; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_13; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_14; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_15; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_32; // @[StoreQueue.scala 75:25:@350.4]
  wire  _GEN_33; // @[StoreQueue.scala 75:25:@350.4]
  wire [3:0] _T_1822; // @[:@372.6]
  wire [3:0] _GEN_35; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_36; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_37; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_38; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_39; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_40; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_41; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_42; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_43; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_44; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_45; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_46; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_47; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_48; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_49; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_66; // @[StoreQueue.scala 75:25:@366.4]
  wire  _GEN_67; // @[StoreQueue.scala 75:25:@366.4]
  wire [3:0] _T_1840; // @[:@388.6]
  wire [3:0] _GEN_69; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_70; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_71; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_72; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_73; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_74; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_75; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_76; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_77; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_78; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_79; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_80; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_81; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_82; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_83; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_100; // @[StoreQueue.scala 75:25:@382.4]
  wire  _GEN_101; // @[StoreQueue.scala 75:25:@382.4]
  wire [3:0] _T_1858; // @[:@404.6]
  wire [3:0] _GEN_103; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_104; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_105; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_106; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_107; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_108; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_109; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_110; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_111; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_112; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_113; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_114; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_115; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_116; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_117; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_134; // @[StoreQueue.scala 75:25:@398.4]
  wire  _GEN_135; // @[StoreQueue.scala 75:25:@398.4]
  wire [3:0] _T_1876; // @[:@420.6]
  wire [3:0] _GEN_137; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_138; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_139; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_140; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_141; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_142; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_143; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_144; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_145; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_146; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_147; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_148; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_149; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_150; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_151; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_168; // @[StoreQueue.scala 75:25:@414.4]
  wire  _GEN_169; // @[StoreQueue.scala 75:25:@414.4]
  wire [3:0] _T_1894; // @[:@436.6]
  wire [3:0] _GEN_171; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_172; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_173; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_174; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_175; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_176; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_177; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_178; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_179; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_180; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_181; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_182; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_183; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_184; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_185; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_202; // @[StoreQueue.scala 75:25:@430.4]
  wire  _GEN_203; // @[StoreQueue.scala 75:25:@430.4]
  wire [3:0] _T_1912; // @[:@452.6]
  wire [3:0] _GEN_205; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_206; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_207; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_208; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_209; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_210; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_211; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_212; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_213; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_214; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_215; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_216; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_217; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_218; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_219; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_236; // @[StoreQueue.scala 75:25:@446.4]
  wire  _GEN_237; // @[StoreQueue.scala 75:25:@446.4]
  wire [3:0] _T_1930; // @[:@468.6]
  wire [3:0] _GEN_239; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_240; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_241; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_242; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_243; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_244; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_245; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_246; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_247; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_248; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_249; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_250; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_251; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_252; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_253; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_270; // @[StoreQueue.scala 75:25:@462.4]
  wire  _GEN_271; // @[StoreQueue.scala 75:25:@462.4]
  wire [3:0] _T_1948; // @[:@484.6]
  wire [3:0] _GEN_273; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_274; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_275; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_276; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_277; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_278; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_279; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_280; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_281; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_282; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_283; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_284; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_285; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_286; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_287; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_304; // @[StoreQueue.scala 75:25:@478.4]
  wire  _GEN_305; // @[StoreQueue.scala 75:25:@478.4]
  wire [3:0] _T_1966; // @[:@500.6]
  wire [3:0] _GEN_307; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_308; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_309; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_310; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_311; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_312; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_313; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_314; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_315; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_316; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_317; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_318; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_319; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_320; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_321; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_338; // @[StoreQueue.scala 75:25:@494.4]
  wire  _GEN_339; // @[StoreQueue.scala 75:25:@494.4]
  wire [3:0] _T_1984; // @[:@516.6]
  wire [3:0] _GEN_341; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_342; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_343; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_344; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_345; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_346; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_347; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_348; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_349; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_350; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_351; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_352; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_353; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_354; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_355; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_372; // @[StoreQueue.scala 75:25:@510.4]
  wire  _GEN_373; // @[StoreQueue.scala 75:25:@510.4]
  wire [3:0] _T_2002; // @[:@532.6]
  wire [3:0] _GEN_375; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_376; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_377; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_378; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_379; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_380; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_381; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_382; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_383; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_384; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_385; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_386; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_387; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_388; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_389; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_406; // @[StoreQueue.scala 75:25:@526.4]
  wire  _GEN_407; // @[StoreQueue.scala 75:25:@526.4]
  wire [3:0] _T_2020; // @[:@548.6]
  wire [3:0] _GEN_409; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_410; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_411; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_412; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_413; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_414; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_415; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_416; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_417; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_418; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_419; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_420; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_421; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_422; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_423; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_440; // @[StoreQueue.scala 75:25:@542.4]
  wire  _GEN_441; // @[StoreQueue.scala 75:25:@542.4]
  wire [3:0] _T_2038; // @[:@564.6]
  wire [3:0] _GEN_443; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_444; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_445; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_446; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_447; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_448; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_449; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_450; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_451; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_452; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_453; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_454; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_455; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_456; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_457; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_474; // @[StoreQueue.scala 75:25:@558.4]
  wire  _GEN_475; // @[StoreQueue.scala 75:25:@558.4]
  wire [3:0] _T_2056; // @[:@580.6]
  wire [3:0] _GEN_477; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_478; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_479; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_480; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_481; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_482; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_483; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_484; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_485; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_486; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_487; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_488; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_489; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_490; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_491; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_508; // @[StoreQueue.scala 75:25:@574.4]
  wire  _GEN_509; // @[StoreQueue.scala 75:25:@574.4]
  wire [3:0] _T_2074; // @[:@596.6]
  wire [3:0] _GEN_511; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_512; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_513; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_514; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_515; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_516; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_517; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_518; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_519; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_520; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_521; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_522; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_523; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_524; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_525; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_542; // @[StoreQueue.scala 75:25:@590.4]
  wire  _GEN_543; // @[StoreQueue.scala 75:25:@590.4]
  reg [3:0] previousLoadHead; // @[StoreQueue.scala 92:33:@606.4]
  reg [31:0] _RAND_146;
  wire [4:0] _T_2096; // @[util.scala 10:8:@615.6]
  wire [4:0] _GEN_31; // @[util.scala 10:14:@616.6]
  wire [4:0] _T_2097; // @[util.scala 10:14:@616.6]
  wire [4:0] _GEN_1203; // @[StoreQueue.scala 96:56:@617.6]
  wire  _T_2098; // @[StoreQueue.scala 96:56:@617.6]
  wire  _T_2099; // @[StoreQueue.scala 95:50:@618.6]
  wire  _T_2101; // @[StoreQueue.scala 95:35:@619.6]
  wire  _T_2103; // @[StoreQueue.scala 100:35:@627.8]
  wire  _T_2104; // @[StoreQueue.scala 100:87:@628.8]
  wire  _T_2105; // @[StoreQueue.scala 100:61:@629.8]
  wire  _T_2107; // @[StoreQueue.scala 102:35:@634.10]
  wire  _T_2108; // @[StoreQueue.scala 103:23:@635.10]
  wire  _T_2109; // @[StoreQueue.scala 103:75:@636.10]
  wire  _T_2110; // @[StoreQueue.scala 103:49:@637.10]
  wire  _T_2112; // @[StoreQueue.scala 103:9:@638.10]
  wire  _T_2113; // @[StoreQueue.scala 102:49:@639.10]
  wire  _GEN_560; // @[StoreQueue.scala 103:96:@640.10]
  wire  _GEN_561; // @[StoreQueue.scala 100:102:@630.8]
  wire  _GEN_562; // @[StoreQueue.scala 98:26:@623.6]
  wire  _GEN_563; // @[StoreQueue.scala 94:35:@608.4]
  wire [4:0] _T_2126; // @[util.scala 10:8:@651.6]
  wire [4:0] _GEN_34; // @[util.scala 10:14:@652.6]
  wire [4:0] _T_2127; // @[util.scala 10:14:@652.6]
  wire  _T_2128; // @[StoreQueue.scala 96:56:@653.6]
  wire  _T_2129; // @[StoreQueue.scala 95:50:@654.6]
  wire  _T_2131; // @[StoreQueue.scala 95:35:@655.6]
  wire  _T_2133; // @[StoreQueue.scala 100:35:@663.8]
  wire  _T_2134; // @[StoreQueue.scala 100:87:@664.8]
  wire  _T_2135; // @[StoreQueue.scala 100:61:@665.8]
  wire  _T_2138; // @[StoreQueue.scala 103:23:@671.10]
  wire  _T_2139; // @[StoreQueue.scala 103:75:@672.10]
  wire  _T_2140; // @[StoreQueue.scala 103:49:@673.10]
  wire  _T_2142; // @[StoreQueue.scala 103:9:@674.10]
  wire  _T_2143; // @[StoreQueue.scala 102:49:@675.10]
  wire  _GEN_580; // @[StoreQueue.scala 103:96:@676.10]
  wire  _GEN_581; // @[StoreQueue.scala 100:102:@666.8]
  wire  _GEN_582; // @[StoreQueue.scala 98:26:@659.6]
  wire  _GEN_583; // @[StoreQueue.scala 94:35:@644.4]
  wire [4:0] _T_2156; // @[util.scala 10:8:@687.6]
  wire [4:0] _GEN_50; // @[util.scala 10:14:@688.6]
  wire [4:0] _T_2157; // @[util.scala 10:14:@688.6]
  wire  _T_2158; // @[StoreQueue.scala 96:56:@689.6]
  wire  _T_2159; // @[StoreQueue.scala 95:50:@690.6]
  wire  _T_2161; // @[StoreQueue.scala 95:35:@691.6]
  wire  _T_2163; // @[StoreQueue.scala 100:35:@699.8]
  wire  _T_2164; // @[StoreQueue.scala 100:87:@700.8]
  wire  _T_2165; // @[StoreQueue.scala 100:61:@701.8]
  wire  _T_2168; // @[StoreQueue.scala 103:23:@707.10]
  wire  _T_2169; // @[StoreQueue.scala 103:75:@708.10]
  wire  _T_2170; // @[StoreQueue.scala 103:49:@709.10]
  wire  _T_2172; // @[StoreQueue.scala 103:9:@710.10]
  wire  _T_2173; // @[StoreQueue.scala 102:49:@711.10]
  wire  _GEN_600; // @[StoreQueue.scala 103:96:@712.10]
  wire  _GEN_601; // @[StoreQueue.scala 100:102:@702.8]
  wire  _GEN_602; // @[StoreQueue.scala 98:26:@695.6]
  wire  _GEN_603; // @[StoreQueue.scala 94:35:@680.4]
  wire [4:0] _T_2186; // @[util.scala 10:8:@723.6]
  wire [4:0] _GEN_51; // @[util.scala 10:14:@724.6]
  wire [4:0] _T_2187; // @[util.scala 10:14:@724.6]
  wire  _T_2188; // @[StoreQueue.scala 96:56:@725.6]
  wire  _T_2189; // @[StoreQueue.scala 95:50:@726.6]
  wire  _T_2191; // @[StoreQueue.scala 95:35:@727.6]
  wire  _T_2193; // @[StoreQueue.scala 100:35:@735.8]
  wire  _T_2194; // @[StoreQueue.scala 100:87:@736.8]
  wire  _T_2195; // @[StoreQueue.scala 100:61:@737.8]
  wire  _T_2198; // @[StoreQueue.scala 103:23:@743.10]
  wire  _T_2199; // @[StoreQueue.scala 103:75:@744.10]
  wire  _T_2200; // @[StoreQueue.scala 103:49:@745.10]
  wire  _T_2202; // @[StoreQueue.scala 103:9:@746.10]
  wire  _T_2203; // @[StoreQueue.scala 102:49:@747.10]
  wire  _GEN_620; // @[StoreQueue.scala 103:96:@748.10]
  wire  _GEN_621; // @[StoreQueue.scala 100:102:@738.8]
  wire  _GEN_622; // @[StoreQueue.scala 98:26:@731.6]
  wire  _GEN_623; // @[StoreQueue.scala 94:35:@716.4]
  wire [4:0] _T_2216; // @[util.scala 10:8:@759.6]
  wire [4:0] _GEN_52; // @[util.scala 10:14:@760.6]
  wire [4:0] _T_2217; // @[util.scala 10:14:@760.6]
  wire  _T_2218; // @[StoreQueue.scala 96:56:@761.6]
  wire  _T_2219; // @[StoreQueue.scala 95:50:@762.6]
  wire  _T_2221; // @[StoreQueue.scala 95:35:@763.6]
  wire  _T_2223; // @[StoreQueue.scala 100:35:@771.8]
  wire  _T_2224; // @[StoreQueue.scala 100:87:@772.8]
  wire  _T_2225; // @[StoreQueue.scala 100:61:@773.8]
  wire  _T_2228; // @[StoreQueue.scala 103:23:@779.10]
  wire  _T_2229; // @[StoreQueue.scala 103:75:@780.10]
  wire  _T_2230; // @[StoreQueue.scala 103:49:@781.10]
  wire  _T_2232; // @[StoreQueue.scala 103:9:@782.10]
  wire  _T_2233; // @[StoreQueue.scala 102:49:@783.10]
  wire  _GEN_640; // @[StoreQueue.scala 103:96:@784.10]
  wire  _GEN_641; // @[StoreQueue.scala 100:102:@774.8]
  wire  _GEN_642; // @[StoreQueue.scala 98:26:@767.6]
  wire  _GEN_643; // @[StoreQueue.scala 94:35:@752.4]
  wire [4:0] _T_2246; // @[util.scala 10:8:@795.6]
  wire [4:0] _GEN_53; // @[util.scala 10:14:@796.6]
  wire [4:0] _T_2247; // @[util.scala 10:14:@796.6]
  wire  _T_2248; // @[StoreQueue.scala 96:56:@797.6]
  wire  _T_2249; // @[StoreQueue.scala 95:50:@798.6]
  wire  _T_2251; // @[StoreQueue.scala 95:35:@799.6]
  wire  _T_2253; // @[StoreQueue.scala 100:35:@807.8]
  wire  _T_2254; // @[StoreQueue.scala 100:87:@808.8]
  wire  _T_2255; // @[StoreQueue.scala 100:61:@809.8]
  wire  _T_2258; // @[StoreQueue.scala 103:23:@815.10]
  wire  _T_2259; // @[StoreQueue.scala 103:75:@816.10]
  wire  _T_2260; // @[StoreQueue.scala 103:49:@817.10]
  wire  _T_2262; // @[StoreQueue.scala 103:9:@818.10]
  wire  _T_2263; // @[StoreQueue.scala 102:49:@819.10]
  wire  _GEN_660; // @[StoreQueue.scala 103:96:@820.10]
  wire  _GEN_661; // @[StoreQueue.scala 100:102:@810.8]
  wire  _GEN_662; // @[StoreQueue.scala 98:26:@803.6]
  wire  _GEN_663; // @[StoreQueue.scala 94:35:@788.4]
  wire [4:0] _T_2276; // @[util.scala 10:8:@831.6]
  wire [4:0] _GEN_54; // @[util.scala 10:14:@832.6]
  wire [4:0] _T_2277; // @[util.scala 10:14:@832.6]
  wire  _T_2278; // @[StoreQueue.scala 96:56:@833.6]
  wire  _T_2279; // @[StoreQueue.scala 95:50:@834.6]
  wire  _T_2281; // @[StoreQueue.scala 95:35:@835.6]
  wire  _T_2283; // @[StoreQueue.scala 100:35:@843.8]
  wire  _T_2284; // @[StoreQueue.scala 100:87:@844.8]
  wire  _T_2285; // @[StoreQueue.scala 100:61:@845.8]
  wire  _T_2288; // @[StoreQueue.scala 103:23:@851.10]
  wire  _T_2289; // @[StoreQueue.scala 103:75:@852.10]
  wire  _T_2290; // @[StoreQueue.scala 103:49:@853.10]
  wire  _T_2292; // @[StoreQueue.scala 103:9:@854.10]
  wire  _T_2293; // @[StoreQueue.scala 102:49:@855.10]
  wire  _GEN_680; // @[StoreQueue.scala 103:96:@856.10]
  wire  _GEN_681; // @[StoreQueue.scala 100:102:@846.8]
  wire  _GEN_682; // @[StoreQueue.scala 98:26:@839.6]
  wire  _GEN_683; // @[StoreQueue.scala 94:35:@824.4]
  wire [4:0] _T_2306; // @[util.scala 10:8:@867.6]
  wire [4:0] _GEN_55; // @[util.scala 10:14:@868.6]
  wire [4:0] _T_2307; // @[util.scala 10:14:@868.6]
  wire  _T_2308; // @[StoreQueue.scala 96:56:@869.6]
  wire  _T_2309; // @[StoreQueue.scala 95:50:@870.6]
  wire  _T_2311; // @[StoreQueue.scala 95:35:@871.6]
  wire  _T_2313; // @[StoreQueue.scala 100:35:@879.8]
  wire  _T_2314; // @[StoreQueue.scala 100:87:@880.8]
  wire  _T_2315; // @[StoreQueue.scala 100:61:@881.8]
  wire  _T_2318; // @[StoreQueue.scala 103:23:@887.10]
  wire  _T_2319; // @[StoreQueue.scala 103:75:@888.10]
  wire  _T_2320; // @[StoreQueue.scala 103:49:@889.10]
  wire  _T_2322; // @[StoreQueue.scala 103:9:@890.10]
  wire  _T_2323; // @[StoreQueue.scala 102:49:@891.10]
  wire  _GEN_700; // @[StoreQueue.scala 103:96:@892.10]
  wire  _GEN_701; // @[StoreQueue.scala 100:102:@882.8]
  wire  _GEN_702; // @[StoreQueue.scala 98:26:@875.6]
  wire  _GEN_703; // @[StoreQueue.scala 94:35:@860.4]
  wire [4:0] _T_2336; // @[util.scala 10:8:@903.6]
  wire [4:0] _GEN_56; // @[util.scala 10:14:@904.6]
  wire [4:0] _T_2337; // @[util.scala 10:14:@904.6]
  wire  _T_2338; // @[StoreQueue.scala 96:56:@905.6]
  wire  _T_2339; // @[StoreQueue.scala 95:50:@906.6]
  wire  _T_2341; // @[StoreQueue.scala 95:35:@907.6]
  wire  _T_2343; // @[StoreQueue.scala 100:35:@915.8]
  wire  _T_2344; // @[StoreQueue.scala 100:87:@916.8]
  wire  _T_2345; // @[StoreQueue.scala 100:61:@917.8]
  wire  _T_2348; // @[StoreQueue.scala 103:23:@923.10]
  wire  _T_2349; // @[StoreQueue.scala 103:75:@924.10]
  wire  _T_2350; // @[StoreQueue.scala 103:49:@925.10]
  wire  _T_2352; // @[StoreQueue.scala 103:9:@926.10]
  wire  _T_2353; // @[StoreQueue.scala 102:49:@927.10]
  wire  _GEN_720; // @[StoreQueue.scala 103:96:@928.10]
  wire  _GEN_721; // @[StoreQueue.scala 100:102:@918.8]
  wire  _GEN_722; // @[StoreQueue.scala 98:26:@911.6]
  wire  _GEN_723; // @[StoreQueue.scala 94:35:@896.4]
  wire [4:0] _T_2366; // @[util.scala 10:8:@939.6]
  wire [4:0] _GEN_57; // @[util.scala 10:14:@940.6]
  wire [4:0] _T_2367; // @[util.scala 10:14:@940.6]
  wire  _T_2368; // @[StoreQueue.scala 96:56:@941.6]
  wire  _T_2369; // @[StoreQueue.scala 95:50:@942.6]
  wire  _T_2371; // @[StoreQueue.scala 95:35:@943.6]
  wire  _T_2373; // @[StoreQueue.scala 100:35:@951.8]
  wire  _T_2374; // @[StoreQueue.scala 100:87:@952.8]
  wire  _T_2375; // @[StoreQueue.scala 100:61:@953.8]
  wire  _T_2378; // @[StoreQueue.scala 103:23:@959.10]
  wire  _T_2379; // @[StoreQueue.scala 103:75:@960.10]
  wire  _T_2380; // @[StoreQueue.scala 103:49:@961.10]
  wire  _T_2382; // @[StoreQueue.scala 103:9:@962.10]
  wire  _T_2383; // @[StoreQueue.scala 102:49:@963.10]
  wire  _GEN_740; // @[StoreQueue.scala 103:96:@964.10]
  wire  _GEN_741; // @[StoreQueue.scala 100:102:@954.8]
  wire  _GEN_742; // @[StoreQueue.scala 98:26:@947.6]
  wire  _GEN_743; // @[StoreQueue.scala 94:35:@932.4]
  wire [4:0] _T_2396; // @[util.scala 10:8:@975.6]
  wire [4:0] _GEN_58; // @[util.scala 10:14:@976.6]
  wire [4:0] _T_2397; // @[util.scala 10:14:@976.6]
  wire  _T_2398; // @[StoreQueue.scala 96:56:@977.6]
  wire  _T_2399; // @[StoreQueue.scala 95:50:@978.6]
  wire  _T_2401; // @[StoreQueue.scala 95:35:@979.6]
  wire  _T_2403; // @[StoreQueue.scala 100:35:@987.8]
  wire  _T_2404; // @[StoreQueue.scala 100:87:@988.8]
  wire  _T_2405; // @[StoreQueue.scala 100:61:@989.8]
  wire  _T_2408; // @[StoreQueue.scala 103:23:@995.10]
  wire  _T_2409; // @[StoreQueue.scala 103:75:@996.10]
  wire  _T_2410; // @[StoreQueue.scala 103:49:@997.10]
  wire  _T_2412; // @[StoreQueue.scala 103:9:@998.10]
  wire  _T_2413; // @[StoreQueue.scala 102:49:@999.10]
  wire  _GEN_760; // @[StoreQueue.scala 103:96:@1000.10]
  wire  _GEN_761; // @[StoreQueue.scala 100:102:@990.8]
  wire  _GEN_762; // @[StoreQueue.scala 98:26:@983.6]
  wire  _GEN_763; // @[StoreQueue.scala 94:35:@968.4]
  wire [4:0] _T_2426; // @[util.scala 10:8:@1011.6]
  wire [4:0] _GEN_59; // @[util.scala 10:14:@1012.6]
  wire [4:0] _T_2427; // @[util.scala 10:14:@1012.6]
  wire  _T_2428; // @[StoreQueue.scala 96:56:@1013.6]
  wire  _T_2429; // @[StoreQueue.scala 95:50:@1014.6]
  wire  _T_2431; // @[StoreQueue.scala 95:35:@1015.6]
  wire  _T_2433; // @[StoreQueue.scala 100:35:@1023.8]
  wire  _T_2434; // @[StoreQueue.scala 100:87:@1024.8]
  wire  _T_2435; // @[StoreQueue.scala 100:61:@1025.8]
  wire  _T_2438; // @[StoreQueue.scala 103:23:@1031.10]
  wire  _T_2439; // @[StoreQueue.scala 103:75:@1032.10]
  wire  _T_2440; // @[StoreQueue.scala 103:49:@1033.10]
  wire  _T_2442; // @[StoreQueue.scala 103:9:@1034.10]
  wire  _T_2443; // @[StoreQueue.scala 102:49:@1035.10]
  wire  _GEN_780; // @[StoreQueue.scala 103:96:@1036.10]
  wire  _GEN_781; // @[StoreQueue.scala 100:102:@1026.8]
  wire  _GEN_782; // @[StoreQueue.scala 98:26:@1019.6]
  wire  _GEN_783; // @[StoreQueue.scala 94:35:@1004.4]
  wire [4:0] _T_2456; // @[util.scala 10:8:@1047.6]
  wire [4:0] _GEN_60; // @[util.scala 10:14:@1048.6]
  wire [4:0] _T_2457; // @[util.scala 10:14:@1048.6]
  wire  _T_2458; // @[StoreQueue.scala 96:56:@1049.6]
  wire  _T_2459; // @[StoreQueue.scala 95:50:@1050.6]
  wire  _T_2461; // @[StoreQueue.scala 95:35:@1051.6]
  wire  _T_2463; // @[StoreQueue.scala 100:35:@1059.8]
  wire  _T_2464; // @[StoreQueue.scala 100:87:@1060.8]
  wire  _T_2465; // @[StoreQueue.scala 100:61:@1061.8]
  wire  _T_2468; // @[StoreQueue.scala 103:23:@1067.10]
  wire  _T_2469; // @[StoreQueue.scala 103:75:@1068.10]
  wire  _T_2470; // @[StoreQueue.scala 103:49:@1069.10]
  wire  _T_2472; // @[StoreQueue.scala 103:9:@1070.10]
  wire  _T_2473; // @[StoreQueue.scala 102:49:@1071.10]
  wire  _GEN_800; // @[StoreQueue.scala 103:96:@1072.10]
  wire  _GEN_801; // @[StoreQueue.scala 100:102:@1062.8]
  wire  _GEN_802; // @[StoreQueue.scala 98:26:@1055.6]
  wire  _GEN_803; // @[StoreQueue.scala 94:35:@1040.4]
  wire [4:0] _T_2486; // @[util.scala 10:8:@1083.6]
  wire [4:0] _GEN_61; // @[util.scala 10:14:@1084.6]
  wire [4:0] _T_2487; // @[util.scala 10:14:@1084.6]
  wire  _T_2488; // @[StoreQueue.scala 96:56:@1085.6]
  wire  _T_2489; // @[StoreQueue.scala 95:50:@1086.6]
  wire  _T_2491; // @[StoreQueue.scala 95:35:@1087.6]
  wire  _T_2493; // @[StoreQueue.scala 100:35:@1095.8]
  wire  _T_2494; // @[StoreQueue.scala 100:87:@1096.8]
  wire  _T_2495; // @[StoreQueue.scala 100:61:@1097.8]
  wire  _T_2498; // @[StoreQueue.scala 103:23:@1103.10]
  wire  _T_2499; // @[StoreQueue.scala 103:75:@1104.10]
  wire  _T_2500; // @[StoreQueue.scala 103:49:@1105.10]
  wire  _T_2502; // @[StoreQueue.scala 103:9:@1106.10]
  wire  _T_2503; // @[StoreQueue.scala 102:49:@1107.10]
  wire  _GEN_820; // @[StoreQueue.scala 103:96:@1108.10]
  wire  _GEN_821; // @[StoreQueue.scala 100:102:@1098.8]
  wire  _GEN_822; // @[StoreQueue.scala 98:26:@1091.6]
  wire  _GEN_823; // @[StoreQueue.scala 94:35:@1076.4]
  wire [4:0] _T_2516; // @[util.scala 10:8:@1119.6]
  wire [4:0] _GEN_62; // @[util.scala 10:14:@1120.6]
  wire [4:0] _T_2517; // @[util.scala 10:14:@1120.6]
  wire  _T_2518; // @[StoreQueue.scala 96:56:@1121.6]
  wire  _T_2519; // @[StoreQueue.scala 95:50:@1122.6]
  wire  _T_2521; // @[StoreQueue.scala 95:35:@1123.6]
  wire  _T_2523; // @[StoreQueue.scala 100:35:@1131.8]
  wire  _T_2524; // @[StoreQueue.scala 100:87:@1132.8]
  wire  _T_2525; // @[StoreQueue.scala 100:61:@1133.8]
  wire  _T_2528; // @[StoreQueue.scala 103:23:@1139.10]
  wire  _T_2529; // @[StoreQueue.scala 103:75:@1140.10]
  wire  _T_2530; // @[StoreQueue.scala 103:49:@1141.10]
  wire  _T_2532; // @[StoreQueue.scala 103:9:@1142.10]
  wire  _T_2533; // @[StoreQueue.scala 102:49:@1143.10]
  wire  _GEN_840; // @[StoreQueue.scala 103:96:@1144.10]
  wire  _GEN_841; // @[StoreQueue.scala 100:102:@1134.8]
  wire  _GEN_842; // @[StoreQueue.scala 98:26:@1127.6]
  wire  _GEN_843; // @[StoreQueue.scala 94:35:@1112.4]
  wire [4:0] _T_2546; // @[util.scala 10:8:@1155.6]
  wire [4:0] _GEN_63; // @[util.scala 10:14:@1156.6]
  wire [4:0] _T_2547; // @[util.scala 10:14:@1156.6]
  wire  _T_2548; // @[StoreQueue.scala 96:56:@1157.6]
  wire  _T_2549; // @[StoreQueue.scala 95:50:@1158.6]
  wire  _T_2551; // @[StoreQueue.scala 95:35:@1159.6]
  wire  _T_2553; // @[StoreQueue.scala 100:35:@1167.8]
  wire  _T_2554; // @[StoreQueue.scala 100:87:@1168.8]
  wire  _T_2555; // @[StoreQueue.scala 100:61:@1169.8]
  wire  _T_2558; // @[StoreQueue.scala 103:23:@1175.10]
  wire  _T_2559; // @[StoreQueue.scala 103:75:@1176.10]
  wire  _T_2560; // @[StoreQueue.scala 103:49:@1177.10]
  wire  _T_2562; // @[StoreQueue.scala 103:9:@1178.10]
  wire  _T_2563; // @[StoreQueue.scala 102:49:@1179.10]
  wire  _GEN_860; // @[StoreQueue.scala 103:96:@1180.10]
  wire  _GEN_861; // @[StoreQueue.scala 100:102:@1170.8]
  wire  _GEN_862; // @[StoreQueue.scala 98:26:@1163.6]
  wire  _GEN_863; // @[StoreQueue.scala 94:35:@1148.4]
  wire  _T_2565; // @[StoreQueue.scala 119:103:@1184.4]
  wire  _T_2567; // @[StoreQueue.scala 120:17:@1185.4]
  wire  _T_2569; // @[StoreQueue.scala 120:35:@1186.4]
  wire  _T_2570; // @[StoreQueue.scala 120:26:@1187.4]
  wire  _T_2572; // @[StoreQueue.scala 120:50:@1188.4]
  wire  _T_2574; // @[StoreQueue.scala 120:81:@1189.4]
  wire  _T_2576; // @[StoreQueue.scala 120:99:@1190.4]
  wire  _T_2577; // @[StoreQueue.scala 120:90:@1191.4]
  wire  _T_2579; // @[StoreQueue.scala 120:67:@1192.4]
  wire  _T_2580; // @[StoreQueue.scala 120:64:@1193.4]
  wire  validEntriesInLoadQ_0; // @[StoreQueue.scala 119:90:@1194.4]
  wire  _T_2584; // @[StoreQueue.scala 120:17:@1196.4]
  wire  _T_2586; // @[StoreQueue.scala 120:35:@1197.4]
  wire  _T_2587; // @[StoreQueue.scala 120:26:@1198.4]
  wire  _T_2591; // @[StoreQueue.scala 120:81:@1200.4]
  wire  _T_2593; // @[StoreQueue.scala 120:99:@1201.4]
  wire  _T_2594; // @[StoreQueue.scala 120:90:@1202.4]
  wire  _T_2596; // @[StoreQueue.scala 120:67:@1203.4]
  wire  _T_2597; // @[StoreQueue.scala 120:64:@1204.4]
  wire  validEntriesInLoadQ_1; // @[StoreQueue.scala 119:90:@1205.4]
  wire  _T_2601; // @[StoreQueue.scala 120:17:@1207.4]
  wire  _T_2603; // @[StoreQueue.scala 120:35:@1208.4]
  wire  _T_2604; // @[StoreQueue.scala 120:26:@1209.4]
  wire  _T_2608; // @[StoreQueue.scala 120:81:@1211.4]
  wire  _T_2610; // @[StoreQueue.scala 120:99:@1212.4]
  wire  _T_2611; // @[StoreQueue.scala 120:90:@1213.4]
  wire  _T_2613; // @[StoreQueue.scala 120:67:@1214.4]
  wire  _T_2614; // @[StoreQueue.scala 120:64:@1215.4]
  wire  validEntriesInLoadQ_2; // @[StoreQueue.scala 119:90:@1216.4]
  wire  _T_2618; // @[StoreQueue.scala 120:17:@1218.4]
  wire  _T_2620; // @[StoreQueue.scala 120:35:@1219.4]
  wire  _T_2621; // @[StoreQueue.scala 120:26:@1220.4]
  wire  _T_2625; // @[StoreQueue.scala 120:81:@1222.4]
  wire  _T_2627; // @[StoreQueue.scala 120:99:@1223.4]
  wire  _T_2628; // @[StoreQueue.scala 120:90:@1224.4]
  wire  _T_2630; // @[StoreQueue.scala 120:67:@1225.4]
  wire  _T_2631; // @[StoreQueue.scala 120:64:@1226.4]
  wire  validEntriesInLoadQ_3; // @[StoreQueue.scala 119:90:@1227.4]
  wire  _T_2635; // @[StoreQueue.scala 120:17:@1229.4]
  wire  _T_2637; // @[StoreQueue.scala 120:35:@1230.4]
  wire  _T_2638; // @[StoreQueue.scala 120:26:@1231.4]
  wire  _T_2642; // @[StoreQueue.scala 120:81:@1233.4]
  wire  _T_2644; // @[StoreQueue.scala 120:99:@1234.4]
  wire  _T_2645; // @[StoreQueue.scala 120:90:@1235.4]
  wire  _T_2647; // @[StoreQueue.scala 120:67:@1236.4]
  wire  _T_2648; // @[StoreQueue.scala 120:64:@1237.4]
  wire  validEntriesInLoadQ_4; // @[StoreQueue.scala 119:90:@1238.4]
  wire  _T_2652; // @[StoreQueue.scala 120:17:@1240.4]
  wire  _T_2654; // @[StoreQueue.scala 120:35:@1241.4]
  wire  _T_2655; // @[StoreQueue.scala 120:26:@1242.4]
  wire  _T_2659; // @[StoreQueue.scala 120:81:@1244.4]
  wire  _T_2661; // @[StoreQueue.scala 120:99:@1245.4]
  wire  _T_2662; // @[StoreQueue.scala 120:90:@1246.4]
  wire  _T_2664; // @[StoreQueue.scala 120:67:@1247.4]
  wire  _T_2665; // @[StoreQueue.scala 120:64:@1248.4]
  wire  validEntriesInLoadQ_5; // @[StoreQueue.scala 119:90:@1249.4]
  wire  _T_2669; // @[StoreQueue.scala 120:17:@1251.4]
  wire  _T_2671; // @[StoreQueue.scala 120:35:@1252.4]
  wire  _T_2672; // @[StoreQueue.scala 120:26:@1253.4]
  wire  _T_2676; // @[StoreQueue.scala 120:81:@1255.4]
  wire  _T_2678; // @[StoreQueue.scala 120:99:@1256.4]
  wire  _T_2679; // @[StoreQueue.scala 120:90:@1257.4]
  wire  _T_2681; // @[StoreQueue.scala 120:67:@1258.4]
  wire  _T_2682; // @[StoreQueue.scala 120:64:@1259.4]
  wire  validEntriesInLoadQ_6; // @[StoreQueue.scala 119:90:@1260.4]
  wire  _T_2686; // @[StoreQueue.scala 120:17:@1262.4]
  wire  _T_2688; // @[StoreQueue.scala 120:35:@1263.4]
  wire  _T_2689; // @[StoreQueue.scala 120:26:@1264.4]
  wire  _T_2693; // @[StoreQueue.scala 120:81:@1266.4]
  wire  _T_2695; // @[StoreQueue.scala 120:99:@1267.4]
  wire  _T_2696; // @[StoreQueue.scala 120:90:@1268.4]
  wire  _T_2698; // @[StoreQueue.scala 120:67:@1269.4]
  wire  _T_2699; // @[StoreQueue.scala 120:64:@1270.4]
  wire  validEntriesInLoadQ_7; // @[StoreQueue.scala 119:90:@1271.4]
  wire  _T_2703; // @[StoreQueue.scala 120:17:@1273.4]
  wire  _T_2705; // @[StoreQueue.scala 120:35:@1274.4]
  wire  _T_2706; // @[StoreQueue.scala 120:26:@1275.4]
  wire  _T_2710; // @[StoreQueue.scala 120:81:@1277.4]
  wire  _T_2712; // @[StoreQueue.scala 120:99:@1278.4]
  wire  _T_2713; // @[StoreQueue.scala 120:90:@1279.4]
  wire  _T_2715; // @[StoreQueue.scala 120:67:@1280.4]
  wire  _T_2716; // @[StoreQueue.scala 120:64:@1281.4]
  wire  validEntriesInLoadQ_8; // @[StoreQueue.scala 119:90:@1282.4]
  wire  _T_2720; // @[StoreQueue.scala 120:17:@1284.4]
  wire  _T_2722; // @[StoreQueue.scala 120:35:@1285.4]
  wire  _T_2723; // @[StoreQueue.scala 120:26:@1286.4]
  wire  _T_2727; // @[StoreQueue.scala 120:81:@1288.4]
  wire  _T_2729; // @[StoreQueue.scala 120:99:@1289.4]
  wire  _T_2730; // @[StoreQueue.scala 120:90:@1290.4]
  wire  _T_2732; // @[StoreQueue.scala 120:67:@1291.4]
  wire  _T_2733; // @[StoreQueue.scala 120:64:@1292.4]
  wire  validEntriesInLoadQ_9; // @[StoreQueue.scala 119:90:@1293.4]
  wire  _T_2737; // @[StoreQueue.scala 120:17:@1295.4]
  wire  _T_2739; // @[StoreQueue.scala 120:35:@1296.4]
  wire  _T_2740; // @[StoreQueue.scala 120:26:@1297.4]
  wire  _T_2744; // @[StoreQueue.scala 120:81:@1299.4]
  wire  _T_2746; // @[StoreQueue.scala 120:99:@1300.4]
  wire  _T_2747; // @[StoreQueue.scala 120:90:@1301.4]
  wire  _T_2749; // @[StoreQueue.scala 120:67:@1302.4]
  wire  _T_2750; // @[StoreQueue.scala 120:64:@1303.4]
  wire  validEntriesInLoadQ_10; // @[StoreQueue.scala 119:90:@1304.4]
  wire  _T_2754; // @[StoreQueue.scala 120:17:@1306.4]
  wire  _T_2756; // @[StoreQueue.scala 120:35:@1307.4]
  wire  _T_2757; // @[StoreQueue.scala 120:26:@1308.4]
  wire  _T_2761; // @[StoreQueue.scala 120:81:@1310.4]
  wire  _T_2763; // @[StoreQueue.scala 120:99:@1311.4]
  wire  _T_2764; // @[StoreQueue.scala 120:90:@1312.4]
  wire  _T_2766; // @[StoreQueue.scala 120:67:@1313.4]
  wire  _T_2767; // @[StoreQueue.scala 120:64:@1314.4]
  wire  validEntriesInLoadQ_11; // @[StoreQueue.scala 119:90:@1315.4]
  wire  _T_2771; // @[StoreQueue.scala 120:17:@1317.4]
  wire  _T_2773; // @[StoreQueue.scala 120:35:@1318.4]
  wire  _T_2774; // @[StoreQueue.scala 120:26:@1319.4]
  wire  _T_2778; // @[StoreQueue.scala 120:81:@1321.4]
  wire  _T_2780; // @[StoreQueue.scala 120:99:@1322.4]
  wire  _T_2781; // @[StoreQueue.scala 120:90:@1323.4]
  wire  _T_2783; // @[StoreQueue.scala 120:67:@1324.4]
  wire  _T_2784; // @[StoreQueue.scala 120:64:@1325.4]
  wire  validEntriesInLoadQ_12; // @[StoreQueue.scala 119:90:@1326.4]
  wire  _T_2788; // @[StoreQueue.scala 120:17:@1328.4]
  wire  _T_2790; // @[StoreQueue.scala 120:35:@1329.4]
  wire  _T_2791; // @[StoreQueue.scala 120:26:@1330.4]
  wire  _T_2795; // @[StoreQueue.scala 120:81:@1332.4]
  wire  _T_2797; // @[StoreQueue.scala 120:99:@1333.4]
  wire  _T_2798; // @[StoreQueue.scala 120:90:@1334.4]
  wire  _T_2800; // @[StoreQueue.scala 120:67:@1335.4]
  wire  _T_2801; // @[StoreQueue.scala 120:64:@1336.4]
  wire  validEntriesInLoadQ_13; // @[StoreQueue.scala 119:90:@1337.4]
  wire  _T_2805; // @[StoreQueue.scala 120:17:@1339.4]
  wire  _T_2807; // @[StoreQueue.scala 120:35:@1340.4]
  wire  _T_2808; // @[StoreQueue.scala 120:26:@1341.4]
  wire  _T_2812; // @[StoreQueue.scala 120:81:@1343.4]
  wire  _T_2814; // @[StoreQueue.scala 120:99:@1344.4]
  wire  _T_2815; // @[StoreQueue.scala 120:90:@1345.4]
  wire  _T_2817; // @[StoreQueue.scala 120:67:@1346.4]
  wire  _T_2818; // @[StoreQueue.scala 120:64:@1347.4]
  wire  validEntriesInLoadQ_14; // @[StoreQueue.scala 119:90:@1348.4]
  wire  validEntriesInLoadQ_15; // @[StoreQueue.scala 119:90:@1359.4]
  wire [3:0] _GEN_865; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_866; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_867; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_868; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_869; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_870; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_871; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_872; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_873; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_874; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_875; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_876; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_877; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_878; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_879; // @[StoreQueue.scala 126:96:@1377.4]
  wire  _T_2861; // @[StoreQueue.scala 126:96:@1377.4]
  wire  loadsToCheck_0; // @[StoreQueue.scala 126:83:@1385.4]
  wire  _T_2891; // @[StoreQueue.scala 127:37:@1388.4]
  wire  _T_2892; // @[StoreQueue.scala 127:28:@1389.4]
  wire  _T_2897; // @[StoreQueue.scala 127:71:@1390.4]
  wire  _T_2900; // @[StoreQueue.scala 127:79:@1392.4]
  wire  _T_2902; // @[StoreQueue.scala 127:55:@1393.4]
  wire  loadsToCheck_1; // @[StoreQueue.scala 126:83:@1394.4]
  wire  _T_2914; // @[StoreQueue.scala 127:37:@1397.4]
  wire  _T_2915; // @[StoreQueue.scala 127:28:@1398.4]
  wire  _T_2920; // @[StoreQueue.scala 127:71:@1399.4]
  wire  _T_2923; // @[StoreQueue.scala 127:79:@1401.4]
  wire  _T_2925; // @[StoreQueue.scala 127:55:@1402.4]
  wire  loadsToCheck_2; // @[StoreQueue.scala 126:83:@1403.4]
  wire  _T_2937; // @[StoreQueue.scala 127:37:@1406.4]
  wire  _T_2938; // @[StoreQueue.scala 127:28:@1407.4]
  wire  _T_2943; // @[StoreQueue.scala 127:71:@1408.4]
  wire  _T_2946; // @[StoreQueue.scala 127:79:@1410.4]
  wire  _T_2948; // @[StoreQueue.scala 127:55:@1411.4]
  wire  loadsToCheck_3; // @[StoreQueue.scala 126:83:@1412.4]
  wire  _T_2960; // @[StoreQueue.scala 127:37:@1415.4]
  wire  _T_2961; // @[StoreQueue.scala 127:28:@1416.4]
  wire  _T_2966; // @[StoreQueue.scala 127:71:@1417.4]
  wire  _T_2969; // @[StoreQueue.scala 127:79:@1419.4]
  wire  _T_2971; // @[StoreQueue.scala 127:55:@1420.4]
  wire  loadsToCheck_4; // @[StoreQueue.scala 126:83:@1421.4]
  wire  _T_2983; // @[StoreQueue.scala 127:37:@1424.4]
  wire  _T_2984; // @[StoreQueue.scala 127:28:@1425.4]
  wire  _T_2989; // @[StoreQueue.scala 127:71:@1426.4]
  wire  _T_2992; // @[StoreQueue.scala 127:79:@1428.4]
  wire  _T_2994; // @[StoreQueue.scala 127:55:@1429.4]
  wire  loadsToCheck_5; // @[StoreQueue.scala 126:83:@1430.4]
  wire  _T_3006; // @[StoreQueue.scala 127:37:@1433.4]
  wire  _T_3007; // @[StoreQueue.scala 127:28:@1434.4]
  wire  _T_3012; // @[StoreQueue.scala 127:71:@1435.4]
  wire  _T_3015; // @[StoreQueue.scala 127:79:@1437.4]
  wire  _T_3017; // @[StoreQueue.scala 127:55:@1438.4]
  wire  loadsToCheck_6; // @[StoreQueue.scala 126:83:@1439.4]
  wire  _T_3029; // @[StoreQueue.scala 127:37:@1442.4]
  wire  _T_3030; // @[StoreQueue.scala 127:28:@1443.4]
  wire  _T_3035; // @[StoreQueue.scala 127:71:@1444.4]
  wire  _T_3038; // @[StoreQueue.scala 127:79:@1446.4]
  wire  _T_3040; // @[StoreQueue.scala 127:55:@1447.4]
  wire  loadsToCheck_7; // @[StoreQueue.scala 126:83:@1448.4]
  wire  _T_3052; // @[StoreQueue.scala 127:37:@1451.4]
  wire  _T_3053; // @[StoreQueue.scala 127:28:@1452.4]
  wire  _T_3058; // @[StoreQueue.scala 127:71:@1453.4]
  wire  _T_3061; // @[StoreQueue.scala 127:79:@1455.4]
  wire  _T_3063; // @[StoreQueue.scala 127:55:@1456.4]
  wire  loadsToCheck_8; // @[StoreQueue.scala 126:83:@1457.4]
  wire  _T_3075; // @[StoreQueue.scala 127:37:@1460.4]
  wire  _T_3076; // @[StoreQueue.scala 127:28:@1461.4]
  wire  _T_3081; // @[StoreQueue.scala 127:71:@1462.4]
  wire  _T_3084; // @[StoreQueue.scala 127:79:@1464.4]
  wire  _T_3086; // @[StoreQueue.scala 127:55:@1465.4]
  wire  loadsToCheck_9; // @[StoreQueue.scala 126:83:@1466.4]
  wire  _T_3098; // @[StoreQueue.scala 127:37:@1469.4]
  wire  _T_3099; // @[StoreQueue.scala 127:28:@1470.4]
  wire  _T_3104; // @[StoreQueue.scala 127:71:@1471.4]
  wire  _T_3107; // @[StoreQueue.scala 127:79:@1473.4]
  wire  _T_3109; // @[StoreQueue.scala 127:55:@1474.4]
  wire  loadsToCheck_10; // @[StoreQueue.scala 126:83:@1475.4]
  wire  _T_3121; // @[StoreQueue.scala 127:37:@1478.4]
  wire  _T_3122; // @[StoreQueue.scala 127:28:@1479.4]
  wire  _T_3127; // @[StoreQueue.scala 127:71:@1480.4]
  wire  _T_3130; // @[StoreQueue.scala 127:79:@1482.4]
  wire  _T_3132; // @[StoreQueue.scala 127:55:@1483.4]
  wire  loadsToCheck_11; // @[StoreQueue.scala 126:83:@1484.4]
  wire  _T_3144; // @[StoreQueue.scala 127:37:@1487.4]
  wire  _T_3145; // @[StoreQueue.scala 127:28:@1488.4]
  wire  _T_3150; // @[StoreQueue.scala 127:71:@1489.4]
  wire  _T_3153; // @[StoreQueue.scala 127:79:@1491.4]
  wire  _T_3155; // @[StoreQueue.scala 127:55:@1492.4]
  wire  loadsToCheck_12; // @[StoreQueue.scala 126:83:@1493.4]
  wire  _T_3167; // @[StoreQueue.scala 127:37:@1496.4]
  wire  _T_3168; // @[StoreQueue.scala 127:28:@1497.4]
  wire  _T_3173; // @[StoreQueue.scala 127:71:@1498.4]
  wire  _T_3176; // @[StoreQueue.scala 127:79:@1500.4]
  wire  _T_3178; // @[StoreQueue.scala 127:55:@1501.4]
  wire  loadsToCheck_13; // @[StoreQueue.scala 126:83:@1502.4]
  wire  _T_3190; // @[StoreQueue.scala 127:37:@1505.4]
  wire  _T_3191; // @[StoreQueue.scala 127:28:@1506.4]
  wire  _T_3196; // @[StoreQueue.scala 127:71:@1507.4]
  wire  _T_3199; // @[StoreQueue.scala 127:79:@1509.4]
  wire  _T_3201; // @[StoreQueue.scala 127:55:@1510.4]
  wire  loadsToCheck_14; // @[StoreQueue.scala 126:83:@1511.4]
  wire  _T_3213; // @[StoreQueue.scala 127:37:@1514.4]
  wire  loadsToCheck_15; // @[StoreQueue.scala 126:83:@1520.4]
  wire  _T_3247; // @[StoreQueue.scala 133:16:@1538.4]
  wire  _GEN_881; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_882; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_883; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_884; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_885; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_886; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_887; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_888; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_889; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_890; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_891; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_892; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_893; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_894; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_895; // @[StoreQueue.scala 133:24:@1539.4]
  wire  entriesToCheck_0; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _T_3252; // @[StoreQueue.scala 133:16:@1540.4]
  wire  entriesToCheck_1; // @[StoreQueue.scala 133:24:@1541.4]
  wire  _T_3257; // @[StoreQueue.scala 133:16:@1542.4]
  wire  entriesToCheck_2; // @[StoreQueue.scala 133:24:@1543.4]
  wire  _T_3262; // @[StoreQueue.scala 133:16:@1544.4]
  wire  entriesToCheck_3; // @[StoreQueue.scala 133:24:@1545.4]
  wire  _T_3267; // @[StoreQueue.scala 133:16:@1546.4]
  wire  entriesToCheck_4; // @[StoreQueue.scala 133:24:@1547.4]
  wire  _T_3272; // @[StoreQueue.scala 133:16:@1548.4]
  wire  entriesToCheck_5; // @[StoreQueue.scala 133:24:@1549.4]
  wire  _T_3277; // @[StoreQueue.scala 133:16:@1550.4]
  wire  entriesToCheck_6; // @[StoreQueue.scala 133:24:@1551.4]
  wire  _T_3282; // @[StoreQueue.scala 133:16:@1552.4]
  wire  entriesToCheck_7; // @[StoreQueue.scala 133:24:@1553.4]
  wire  _T_3287; // @[StoreQueue.scala 133:16:@1554.4]
  wire  entriesToCheck_8; // @[StoreQueue.scala 133:24:@1555.4]
  wire  _T_3292; // @[StoreQueue.scala 133:16:@1556.4]
  wire  entriesToCheck_9; // @[StoreQueue.scala 133:24:@1557.4]
  wire  _T_3297; // @[StoreQueue.scala 133:16:@1558.4]
  wire  entriesToCheck_10; // @[StoreQueue.scala 133:24:@1559.4]
  wire  _T_3302; // @[StoreQueue.scala 133:16:@1560.4]
  wire  entriesToCheck_11; // @[StoreQueue.scala 133:24:@1561.4]
  wire  _T_3307; // @[StoreQueue.scala 133:16:@1562.4]
  wire  entriesToCheck_12; // @[StoreQueue.scala 133:24:@1563.4]
  wire  _T_3312; // @[StoreQueue.scala 133:16:@1564.4]
  wire  entriesToCheck_13; // @[StoreQueue.scala 133:24:@1565.4]
  wire  _T_3317; // @[StoreQueue.scala 133:16:@1566.4]
  wire  entriesToCheck_14; // @[StoreQueue.scala 133:24:@1567.4]
  wire  _T_3322; // @[StoreQueue.scala 133:16:@1568.4]
  wire  entriesToCheck_15; // @[StoreQueue.scala 133:24:@1569.4]
  wire  _T_3370; // @[StoreQueue.scala 140:34:@1588.4]
  wire  _T_3371; // @[StoreQueue.scala 140:64:@1589.4]
  wire [31:0] _GEN_897; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_898; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_899; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_900; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_901; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_902; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_903; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_904; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_905; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_906; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_907; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_908; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_909; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_910; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_911; // @[StoreQueue.scala 141:51:@1590.4]
  wire  _T_3375; // @[StoreQueue.scala 141:51:@1590.4]
  wire  _T_3376; // @[StoreQueue.scala 141:36:@1591.4]
  wire  noConflicts_0; // @[StoreQueue.scala 140:95:@1592.4]
  wire  _T_3379; // @[StoreQueue.scala 140:34:@1594.4]
  wire  _T_3380; // @[StoreQueue.scala 140:64:@1595.4]
  wire  _T_3384; // @[StoreQueue.scala 141:51:@1596.4]
  wire  _T_3385; // @[StoreQueue.scala 141:36:@1597.4]
  wire  noConflicts_1; // @[StoreQueue.scala 140:95:@1598.4]
  wire  _T_3388; // @[StoreQueue.scala 140:34:@1600.4]
  wire  _T_3389; // @[StoreQueue.scala 140:64:@1601.4]
  wire  _T_3393; // @[StoreQueue.scala 141:51:@1602.4]
  wire  _T_3394; // @[StoreQueue.scala 141:36:@1603.4]
  wire  noConflicts_2; // @[StoreQueue.scala 140:95:@1604.4]
  wire  _T_3397; // @[StoreQueue.scala 140:34:@1606.4]
  wire  _T_3398; // @[StoreQueue.scala 140:64:@1607.4]
  wire  _T_3402; // @[StoreQueue.scala 141:51:@1608.4]
  wire  _T_3403; // @[StoreQueue.scala 141:36:@1609.4]
  wire  noConflicts_3; // @[StoreQueue.scala 140:95:@1610.4]
  wire  _T_3406; // @[StoreQueue.scala 140:34:@1612.4]
  wire  _T_3407; // @[StoreQueue.scala 140:64:@1613.4]
  wire  _T_3411; // @[StoreQueue.scala 141:51:@1614.4]
  wire  _T_3412; // @[StoreQueue.scala 141:36:@1615.4]
  wire  noConflicts_4; // @[StoreQueue.scala 140:95:@1616.4]
  wire  _T_3415; // @[StoreQueue.scala 140:34:@1618.4]
  wire  _T_3416; // @[StoreQueue.scala 140:64:@1619.4]
  wire  _T_3420; // @[StoreQueue.scala 141:51:@1620.4]
  wire  _T_3421; // @[StoreQueue.scala 141:36:@1621.4]
  wire  noConflicts_5; // @[StoreQueue.scala 140:95:@1622.4]
  wire  _T_3424; // @[StoreQueue.scala 140:34:@1624.4]
  wire  _T_3425; // @[StoreQueue.scala 140:64:@1625.4]
  wire  _T_3429; // @[StoreQueue.scala 141:51:@1626.4]
  wire  _T_3430; // @[StoreQueue.scala 141:36:@1627.4]
  wire  noConflicts_6; // @[StoreQueue.scala 140:95:@1628.4]
  wire  _T_3433; // @[StoreQueue.scala 140:34:@1630.4]
  wire  _T_3434; // @[StoreQueue.scala 140:64:@1631.4]
  wire  _T_3438; // @[StoreQueue.scala 141:51:@1632.4]
  wire  _T_3439; // @[StoreQueue.scala 141:36:@1633.4]
  wire  noConflicts_7; // @[StoreQueue.scala 140:95:@1634.4]
  wire  _T_3442; // @[StoreQueue.scala 140:34:@1636.4]
  wire  _T_3443; // @[StoreQueue.scala 140:64:@1637.4]
  wire  _T_3447; // @[StoreQueue.scala 141:51:@1638.4]
  wire  _T_3448; // @[StoreQueue.scala 141:36:@1639.4]
  wire  noConflicts_8; // @[StoreQueue.scala 140:95:@1640.4]
  wire  _T_3451; // @[StoreQueue.scala 140:34:@1642.4]
  wire  _T_3452; // @[StoreQueue.scala 140:64:@1643.4]
  wire  _T_3456; // @[StoreQueue.scala 141:51:@1644.4]
  wire  _T_3457; // @[StoreQueue.scala 141:36:@1645.4]
  wire  noConflicts_9; // @[StoreQueue.scala 140:95:@1646.4]
  wire  _T_3460; // @[StoreQueue.scala 140:34:@1648.4]
  wire  _T_3461; // @[StoreQueue.scala 140:64:@1649.4]
  wire  _T_3465; // @[StoreQueue.scala 141:51:@1650.4]
  wire  _T_3466; // @[StoreQueue.scala 141:36:@1651.4]
  wire  noConflicts_10; // @[StoreQueue.scala 140:95:@1652.4]
  wire  _T_3469; // @[StoreQueue.scala 140:34:@1654.4]
  wire  _T_3470; // @[StoreQueue.scala 140:64:@1655.4]
  wire  _T_3474; // @[StoreQueue.scala 141:51:@1656.4]
  wire  _T_3475; // @[StoreQueue.scala 141:36:@1657.4]
  wire  noConflicts_11; // @[StoreQueue.scala 140:95:@1658.4]
  wire  _T_3478; // @[StoreQueue.scala 140:34:@1660.4]
  wire  _T_3479; // @[StoreQueue.scala 140:64:@1661.4]
  wire  _T_3483; // @[StoreQueue.scala 141:51:@1662.4]
  wire  _T_3484; // @[StoreQueue.scala 141:36:@1663.4]
  wire  noConflicts_12; // @[StoreQueue.scala 140:95:@1664.4]
  wire  _T_3487; // @[StoreQueue.scala 140:34:@1666.4]
  wire  _T_3488; // @[StoreQueue.scala 140:64:@1667.4]
  wire  _T_3492; // @[StoreQueue.scala 141:51:@1668.4]
  wire  _T_3493; // @[StoreQueue.scala 141:36:@1669.4]
  wire  noConflicts_13; // @[StoreQueue.scala 140:95:@1670.4]
  wire  _T_3496; // @[StoreQueue.scala 140:34:@1672.4]
  wire  _T_3497; // @[StoreQueue.scala 140:64:@1673.4]
  wire  _T_3501; // @[StoreQueue.scala 141:51:@1674.4]
  wire  _T_3502; // @[StoreQueue.scala 141:36:@1675.4]
  wire  noConflicts_14; // @[StoreQueue.scala 140:95:@1676.4]
  wire  _T_3505; // @[StoreQueue.scala 140:34:@1678.4]
  wire  _T_3506; // @[StoreQueue.scala 140:64:@1679.4]
  wire  _T_3510; // @[StoreQueue.scala 141:51:@1680.4]
  wire  _T_3511; // @[StoreQueue.scala 141:36:@1681.4]
  wire  noConflicts_15; // @[StoreQueue.scala 140:95:@1682.4]
  wire  _GEN_913; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_914; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_915; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_916; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_917; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_918; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_919; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_920; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_921; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_922; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_923; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_924; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_925; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_926; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_927; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_929; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_930; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_931; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_932; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_933; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_934; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_935; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_936; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_937; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_938; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_939; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_940; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_941; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_942; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_943; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _T_3519; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_945; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_946; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_947; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_948; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_949; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_950; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_951; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_952; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_953; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_954; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_955; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_956; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_957; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_958; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_959; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _T_3524; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _T_3525; // @[StoreQueue.scala 154:63:@1686.4]
  wire  _T_3528; // @[StoreQueue.scala 154:109:@1688.4]
  wire  _T_3529; // @[StoreQueue.scala 154:109:@1689.4]
  wire  _T_3530; // @[StoreQueue.scala 154:109:@1690.4]
  wire  _T_3531; // @[StoreQueue.scala 154:109:@1691.4]
  wire  _T_3532; // @[StoreQueue.scala 154:109:@1692.4]
  wire  _T_3533; // @[StoreQueue.scala 154:109:@1693.4]
  wire  _T_3534; // @[StoreQueue.scala 154:109:@1694.4]
  wire  _T_3535; // @[StoreQueue.scala 154:109:@1695.4]
  wire  _T_3536; // @[StoreQueue.scala 154:109:@1696.4]
  wire  _T_3537; // @[StoreQueue.scala 154:109:@1697.4]
  wire  _T_3538; // @[StoreQueue.scala 154:109:@1698.4]
  wire  _T_3539; // @[StoreQueue.scala 154:109:@1699.4]
  wire  _T_3540; // @[StoreQueue.scala 154:109:@1700.4]
  wire  _T_3541; // @[StoreQueue.scala 154:109:@1701.4]
  wire  _T_3542; // @[StoreQueue.scala 154:109:@1702.4]
  wire  storeRequest; // @[StoreQueue.scala 154:88:@1703.4]
  wire  _T_3545; // @[StoreQueue.scala 164:23:@1708.6]
  wire  _T_3546; // @[StoreQueue.scala 164:43:@1709.6]
  wire  _T_3547; // @[StoreQueue.scala 164:59:@1710.6]
  wire  _GEN_960; // @[StoreQueue.scala 164:86:@1711.6]
  wire  _GEN_961; // @[StoreQueue.scala 162:37:@1704.4]
  wire  _T_3551; // @[StoreQueue.scala 164:23:@1718.6]
  wire  _T_3552; // @[StoreQueue.scala 164:43:@1719.6]
  wire  _T_3553; // @[StoreQueue.scala 164:59:@1720.6]
  wire  _GEN_962; // @[StoreQueue.scala 164:86:@1721.6]
  wire  _GEN_963; // @[StoreQueue.scala 162:37:@1714.4]
  wire  _T_3557; // @[StoreQueue.scala 164:23:@1728.6]
  wire  _T_3558; // @[StoreQueue.scala 164:43:@1729.6]
  wire  _T_3559; // @[StoreQueue.scala 164:59:@1730.6]
  wire  _GEN_964; // @[StoreQueue.scala 164:86:@1731.6]
  wire  _GEN_965; // @[StoreQueue.scala 162:37:@1724.4]
  wire  _T_3563; // @[StoreQueue.scala 164:23:@1738.6]
  wire  _T_3564; // @[StoreQueue.scala 164:43:@1739.6]
  wire  _T_3565; // @[StoreQueue.scala 164:59:@1740.6]
  wire  _GEN_966; // @[StoreQueue.scala 164:86:@1741.6]
  wire  _GEN_967; // @[StoreQueue.scala 162:37:@1734.4]
  wire  _T_3569; // @[StoreQueue.scala 164:23:@1748.6]
  wire  _T_3570; // @[StoreQueue.scala 164:43:@1749.6]
  wire  _T_3571; // @[StoreQueue.scala 164:59:@1750.6]
  wire  _GEN_968; // @[StoreQueue.scala 164:86:@1751.6]
  wire  _GEN_969; // @[StoreQueue.scala 162:37:@1744.4]
  wire  _T_3575; // @[StoreQueue.scala 164:23:@1758.6]
  wire  _T_3576; // @[StoreQueue.scala 164:43:@1759.6]
  wire  _T_3577; // @[StoreQueue.scala 164:59:@1760.6]
  wire  _GEN_970; // @[StoreQueue.scala 164:86:@1761.6]
  wire  _GEN_971; // @[StoreQueue.scala 162:37:@1754.4]
  wire  _T_3581; // @[StoreQueue.scala 164:23:@1768.6]
  wire  _T_3582; // @[StoreQueue.scala 164:43:@1769.6]
  wire  _T_3583; // @[StoreQueue.scala 164:59:@1770.6]
  wire  _GEN_972; // @[StoreQueue.scala 164:86:@1771.6]
  wire  _GEN_973; // @[StoreQueue.scala 162:37:@1764.4]
  wire  _T_3587; // @[StoreQueue.scala 164:23:@1778.6]
  wire  _T_3588; // @[StoreQueue.scala 164:43:@1779.6]
  wire  _T_3589; // @[StoreQueue.scala 164:59:@1780.6]
  wire  _GEN_974; // @[StoreQueue.scala 164:86:@1781.6]
  wire  _GEN_975; // @[StoreQueue.scala 162:37:@1774.4]
  wire  _T_3593; // @[StoreQueue.scala 164:23:@1788.6]
  wire  _T_3594; // @[StoreQueue.scala 164:43:@1789.6]
  wire  _T_3595; // @[StoreQueue.scala 164:59:@1790.6]
  wire  _GEN_976; // @[StoreQueue.scala 164:86:@1791.6]
  wire  _GEN_977; // @[StoreQueue.scala 162:37:@1784.4]
  wire  _T_3599; // @[StoreQueue.scala 164:23:@1798.6]
  wire  _T_3600; // @[StoreQueue.scala 164:43:@1799.6]
  wire  _T_3601; // @[StoreQueue.scala 164:59:@1800.6]
  wire  _GEN_978; // @[StoreQueue.scala 164:86:@1801.6]
  wire  _GEN_979; // @[StoreQueue.scala 162:37:@1794.4]
  wire  _T_3605; // @[StoreQueue.scala 164:23:@1808.6]
  wire  _T_3606; // @[StoreQueue.scala 164:43:@1809.6]
  wire  _T_3607; // @[StoreQueue.scala 164:59:@1810.6]
  wire  _GEN_980; // @[StoreQueue.scala 164:86:@1811.6]
  wire  _GEN_981; // @[StoreQueue.scala 162:37:@1804.4]
  wire  _T_3611; // @[StoreQueue.scala 164:23:@1818.6]
  wire  _T_3612; // @[StoreQueue.scala 164:43:@1819.6]
  wire  _T_3613; // @[StoreQueue.scala 164:59:@1820.6]
  wire  _GEN_982; // @[StoreQueue.scala 164:86:@1821.6]
  wire  _GEN_983; // @[StoreQueue.scala 162:37:@1814.4]
  wire  _T_3617; // @[StoreQueue.scala 164:23:@1828.6]
  wire  _T_3618; // @[StoreQueue.scala 164:43:@1829.6]
  wire  _T_3619; // @[StoreQueue.scala 164:59:@1830.6]
  wire  _GEN_984; // @[StoreQueue.scala 164:86:@1831.6]
  wire  _GEN_985; // @[StoreQueue.scala 162:37:@1824.4]
  wire  _T_3623; // @[StoreQueue.scala 164:23:@1838.6]
  wire  _T_3624; // @[StoreQueue.scala 164:43:@1839.6]
  wire  _T_3625; // @[StoreQueue.scala 164:59:@1840.6]
  wire  _GEN_986; // @[StoreQueue.scala 164:86:@1841.6]
  wire  _GEN_987; // @[StoreQueue.scala 162:37:@1834.4]
  wire  _T_3629; // @[StoreQueue.scala 164:23:@1848.6]
  wire  _T_3630; // @[StoreQueue.scala 164:43:@1849.6]
  wire  _T_3631; // @[StoreQueue.scala 164:59:@1850.6]
  wire  _GEN_988; // @[StoreQueue.scala 164:86:@1851.6]
  wire  _GEN_989; // @[StoreQueue.scala 162:37:@1844.4]
  wire  _T_3635; // @[StoreQueue.scala 164:23:@1858.6]
  wire  _T_3636; // @[StoreQueue.scala 164:43:@1859.6]
  wire  _T_3637; // @[StoreQueue.scala 164:59:@1860.6]
  wire  _GEN_990; // @[StoreQueue.scala 164:86:@1861.6]
  wire  _GEN_991; // @[StoreQueue.scala 162:37:@1854.4]
  wire  entriesPorts_0_0; // @[StoreQueue.scala 180:72:@1865.4]
  wire  entriesPorts_0_1; // @[StoreQueue.scala 180:72:@1867.4]
  wire  entriesPorts_0_2; // @[StoreQueue.scala 180:72:@1869.4]
  wire  entriesPorts_0_3; // @[StoreQueue.scala 180:72:@1871.4]
  wire  entriesPorts_0_4; // @[StoreQueue.scala 180:72:@1873.4]
  wire  entriesPorts_0_5; // @[StoreQueue.scala 180:72:@1875.4]
  wire  entriesPorts_0_6; // @[StoreQueue.scala 180:72:@1877.4]
  wire  entriesPorts_0_7; // @[StoreQueue.scala 180:72:@1879.4]
  wire  entriesPorts_0_8; // @[StoreQueue.scala 180:72:@1881.4]
  wire  entriesPorts_0_9; // @[StoreQueue.scala 180:72:@1883.4]
  wire  entriesPorts_0_10; // @[StoreQueue.scala 180:72:@1885.4]
  wire  entriesPorts_0_11; // @[StoreQueue.scala 180:72:@1887.4]
  wire  entriesPorts_0_12; // @[StoreQueue.scala 180:72:@1889.4]
  wire  entriesPorts_0_13; // @[StoreQueue.scala 180:72:@1891.4]
  wire  entriesPorts_0_14; // @[StoreQueue.scala 180:72:@1893.4]
  wire  entriesPorts_0_15; // @[StoreQueue.scala 180:72:@1895.4]
  wire  _T_4122; // @[StoreQueue.scala 192:91:@1899.4]
  wire  _T_4123; // @[StoreQueue.scala 192:88:@1900.4]
  wire  _T_4125; // @[StoreQueue.scala 192:91:@1901.4]
  wire  _T_4126; // @[StoreQueue.scala 192:88:@1902.4]
  wire  _T_4128; // @[StoreQueue.scala 192:91:@1903.4]
  wire  _T_4129; // @[StoreQueue.scala 192:88:@1904.4]
  wire  _T_4131; // @[StoreQueue.scala 192:91:@1905.4]
  wire  _T_4132; // @[StoreQueue.scala 192:88:@1906.4]
  wire  _T_4134; // @[StoreQueue.scala 192:91:@1907.4]
  wire  _T_4135; // @[StoreQueue.scala 192:88:@1908.4]
  wire  _T_4137; // @[StoreQueue.scala 192:91:@1909.4]
  wire  _T_4138; // @[StoreQueue.scala 192:88:@1910.4]
  wire  _T_4140; // @[StoreQueue.scala 192:91:@1911.4]
  wire  _T_4141; // @[StoreQueue.scala 192:88:@1912.4]
  wire  _T_4143; // @[StoreQueue.scala 192:91:@1913.4]
  wire  _T_4144; // @[StoreQueue.scala 192:88:@1914.4]
  wire  _T_4146; // @[StoreQueue.scala 192:91:@1915.4]
  wire  _T_4147; // @[StoreQueue.scala 192:88:@1916.4]
  wire  _T_4149; // @[StoreQueue.scala 192:91:@1917.4]
  wire  _T_4150; // @[StoreQueue.scala 192:88:@1918.4]
  wire  _T_4152; // @[StoreQueue.scala 192:91:@1919.4]
  wire  _T_4153; // @[StoreQueue.scala 192:88:@1920.4]
  wire  _T_4155; // @[StoreQueue.scala 192:91:@1921.4]
  wire  _T_4156; // @[StoreQueue.scala 192:88:@1922.4]
  wire  _T_4158; // @[StoreQueue.scala 192:91:@1923.4]
  wire  _T_4159; // @[StoreQueue.scala 192:88:@1924.4]
  wire  _T_4161; // @[StoreQueue.scala 192:91:@1925.4]
  wire  _T_4162; // @[StoreQueue.scala 192:88:@1926.4]
  wire  _T_4164; // @[StoreQueue.scala 192:91:@1927.4]
  wire  _T_4165; // @[StoreQueue.scala 192:88:@1928.4]
  wire  _T_4167; // @[StoreQueue.scala 192:91:@1929.4]
  wire  _T_4168; // @[StoreQueue.scala 192:88:@1930.4]
  wire  _T_4192; // @[StoreQueue.scala 193:91:@1948.4]
  wire  _T_4193; // @[StoreQueue.scala 193:88:@1949.4]
  wire  _T_4195; // @[StoreQueue.scala 193:91:@1950.4]
  wire  _T_4196; // @[StoreQueue.scala 193:88:@1951.4]
  wire  _T_4198; // @[StoreQueue.scala 193:91:@1952.4]
  wire  _T_4199; // @[StoreQueue.scala 193:88:@1953.4]
  wire  _T_4201; // @[StoreQueue.scala 193:91:@1954.4]
  wire  _T_4202; // @[StoreQueue.scala 193:88:@1955.4]
  wire  _T_4204; // @[StoreQueue.scala 193:91:@1956.4]
  wire  _T_4205; // @[StoreQueue.scala 193:88:@1957.4]
  wire  _T_4207; // @[StoreQueue.scala 193:91:@1958.4]
  wire  _T_4208; // @[StoreQueue.scala 193:88:@1959.4]
  wire  _T_4210; // @[StoreQueue.scala 193:91:@1960.4]
  wire  _T_4211; // @[StoreQueue.scala 193:88:@1961.4]
  wire  _T_4213; // @[StoreQueue.scala 193:91:@1962.4]
  wire  _T_4214; // @[StoreQueue.scala 193:88:@1963.4]
  wire  _T_4216; // @[StoreQueue.scala 193:91:@1964.4]
  wire  _T_4217; // @[StoreQueue.scala 193:88:@1965.4]
  wire  _T_4219; // @[StoreQueue.scala 193:91:@1966.4]
  wire  _T_4220; // @[StoreQueue.scala 193:88:@1967.4]
  wire  _T_4222; // @[StoreQueue.scala 193:91:@1968.4]
  wire  _T_4223; // @[StoreQueue.scala 193:88:@1969.4]
  wire  _T_4225; // @[StoreQueue.scala 193:91:@1970.4]
  wire  _T_4226; // @[StoreQueue.scala 193:88:@1971.4]
  wire  _T_4228; // @[StoreQueue.scala 193:91:@1972.4]
  wire  _T_4229; // @[StoreQueue.scala 193:88:@1973.4]
  wire  _T_4231; // @[StoreQueue.scala 193:91:@1974.4]
  wire  _T_4232; // @[StoreQueue.scala 193:88:@1975.4]
  wire  _T_4234; // @[StoreQueue.scala 193:91:@1976.4]
  wire  _T_4235; // @[StoreQueue.scala 193:88:@1977.4]
  wire  _T_4237; // @[StoreQueue.scala 193:91:@1978.4]
  wire  _T_4238; // @[StoreQueue.scala 193:88:@1979.4]
  wire [15:0] _T_4263; // @[OneHot.scala 52:12:@1998.4]
  wire  _T_4265; // @[util.scala 33:60:@2000.4]
  wire  _T_4266; // @[util.scala 33:60:@2001.4]
  wire  _T_4267; // @[util.scala 33:60:@2002.4]
  wire  _T_4268; // @[util.scala 33:60:@2003.4]
  wire  _T_4269; // @[util.scala 33:60:@2004.4]
  wire  _T_4270; // @[util.scala 33:60:@2005.4]
  wire  _T_4271; // @[util.scala 33:60:@2006.4]
  wire  _T_4272; // @[util.scala 33:60:@2007.4]
  wire  _T_4273; // @[util.scala 33:60:@2008.4]
  wire  _T_4274; // @[util.scala 33:60:@2009.4]
  wire  _T_4275; // @[util.scala 33:60:@2010.4]
  wire  _T_4276; // @[util.scala 33:60:@2011.4]
  wire  _T_4277; // @[util.scala 33:60:@2012.4]
  wire  _T_4278; // @[util.scala 33:60:@2013.4]
  wire  _T_4279; // @[util.scala 33:60:@2014.4]
  wire  _T_4280; // @[util.scala 33:60:@2015.4]
  wire [15:0] _T_4321; // @[Mux.scala 31:69:@2033.4]
  wire [15:0] _T_4322; // @[Mux.scala 31:69:@2034.4]
  wire [15:0] _T_4323; // @[Mux.scala 31:69:@2035.4]
  wire [15:0] _T_4324; // @[Mux.scala 31:69:@2036.4]
  wire [15:0] _T_4325; // @[Mux.scala 31:69:@2037.4]
  wire [15:0] _T_4326; // @[Mux.scala 31:69:@2038.4]
  wire [15:0] _T_4327; // @[Mux.scala 31:69:@2039.4]
  wire [15:0] _T_4328; // @[Mux.scala 31:69:@2040.4]
  wire [15:0] _T_4329; // @[Mux.scala 31:69:@2041.4]
  wire [15:0] _T_4330; // @[Mux.scala 31:69:@2042.4]
  wire [15:0] _T_4331; // @[Mux.scala 31:69:@2043.4]
  wire [15:0] _T_4332; // @[Mux.scala 31:69:@2044.4]
  wire [15:0] _T_4333; // @[Mux.scala 31:69:@2045.4]
  wire [15:0] _T_4334; // @[Mux.scala 31:69:@2046.4]
  wire [15:0] _T_4335; // @[Mux.scala 31:69:@2047.4]
  wire [15:0] _T_4336; // @[Mux.scala 31:69:@2048.4]
  wire  _T_4337; // @[OneHot.scala 66:30:@2049.4]
  wire  _T_4338; // @[OneHot.scala 66:30:@2050.4]
  wire  _T_4339; // @[OneHot.scala 66:30:@2051.4]
  wire  _T_4340; // @[OneHot.scala 66:30:@2052.4]
  wire  _T_4341; // @[OneHot.scala 66:30:@2053.4]
  wire  _T_4342; // @[OneHot.scala 66:30:@2054.4]
  wire  _T_4343; // @[OneHot.scala 66:30:@2055.4]
  wire  _T_4344; // @[OneHot.scala 66:30:@2056.4]
  wire  _T_4345; // @[OneHot.scala 66:30:@2057.4]
  wire  _T_4346; // @[OneHot.scala 66:30:@2058.4]
  wire  _T_4347; // @[OneHot.scala 66:30:@2059.4]
  wire  _T_4348; // @[OneHot.scala 66:30:@2060.4]
  wire  _T_4349; // @[OneHot.scala 66:30:@2061.4]
  wire  _T_4350; // @[OneHot.scala 66:30:@2062.4]
  wire  _T_4351; // @[OneHot.scala 66:30:@2063.4]
  wire  _T_4352; // @[OneHot.scala 66:30:@2064.4]
  wire [15:0] _T_4393; // @[Mux.scala 31:69:@2082.4]
  wire [15:0] _T_4394; // @[Mux.scala 31:69:@2083.4]
  wire [15:0] _T_4395; // @[Mux.scala 31:69:@2084.4]
  wire [15:0] _T_4396; // @[Mux.scala 31:69:@2085.4]
  wire [15:0] _T_4397; // @[Mux.scala 31:69:@2086.4]
  wire [15:0] _T_4398; // @[Mux.scala 31:69:@2087.4]
  wire [15:0] _T_4399; // @[Mux.scala 31:69:@2088.4]
  wire [15:0] _T_4400; // @[Mux.scala 31:69:@2089.4]
  wire [15:0] _T_4401; // @[Mux.scala 31:69:@2090.4]
  wire [15:0] _T_4402; // @[Mux.scala 31:69:@2091.4]
  wire [15:0] _T_4403; // @[Mux.scala 31:69:@2092.4]
  wire [15:0] _T_4404; // @[Mux.scala 31:69:@2093.4]
  wire [15:0] _T_4405; // @[Mux.scala 31:69:@2094.4]
  wire [15:0] _T_4406; // @[Mux.scala 31:69:@2095.4]
  wire [15:0] _T_4407; // @[Mux.scala 31:69:@2096.4]
  wire [15:0] _T_4408; // @[Mux.scala 31:69:@2097.4]
  wire  _T_4409; // @[OneHot.scala 66:30:@2098.4]
  wire  _T_4410; // @[OneHot.scala 66:30:@2099.4]
  wire  _T_4411; // @[OneHot.scala 66:30:@2100.4]
  wire  _T_4412; // @[OneHot.scala 66:30:@2101.4]
  wire  _T_4413; // @[OneHot.scala 66:30:@2102.4]
  wire  _T_4414; // @[OneHot.scala 66:30:@2103.4]
  wire  _T_4415; // @[OneHot.scala 66:30:@2104.4]
  wire  _T_4416; // @[OneHot.scala 66:30:@2105.4]
  wire  _T_4417; // @[OneHot.scala 66:30:@2106.4]
  wire  _T_4418; // @[OneHot.scala 66:30:@2107.4]
  wire  _T_4419; // @[OneHot.scala 66:30:@2108.4]
  wire  _T_4420; // @[OneHot.scala 66:30:@2109.4]
  wire  _T_4421; // @[OneHot.scala 66:30:@2110.4]
  wire  _T_4422; // @[OneHot.scala 66:30:@2111.4]
  wire  _T_4423; // @[OneHot.scala 66:30:@2112.4]
  wire  _T_4424; // @[OneHot.scala 66:30:@2113.4]
  wire [15:0] _T_4465; // @[Mux.scala 31:69:@2131.4]
  wire [15:0] _T_4466; // @[Mux.scala 31:69:@2132.4]
  wire [15:0] _T_4467; // @[Mux.scala 31:69:@2133.4]
  wire [15:0] _T_4468; // @[Mux.scala 31:69:@2134.4]
  wire [15:0] _T_4469; // @[Mux.scala 31:69:@2135.4]
  wire [15:0] _T_4470; // @[Mux.scala 31:69:@2136.4]
  wire [15:0] _T_4471; // @[Mux.scala 31:69:@2137.4]
  wire [15:0] _T_4472; // @[Mux.scala 31:69:@2138.4]
  wire [15:0] _T_4473; // @[Mux.scala 31:69:@2139.4]
  wire [15:0] _T_4474; // @[Mux.scala 31:69:@2140.4]
  wire [15:0] _T_4475; // @[Mux.scala 31:69:@2141.4]
  wire [15:0] _T_4476; // @[Mux.scala 31:69:@2142.4]
  wire [15:0] _T_4477; // @[Mux.scala 31:69:@2143.4]
  wire [15:0] _T_4478; // @[Mux.scala 31:69:@2144.4]
  wire [15:0] _T_4479; // @[Mux.scala 31:69:@2145.4]
  wire [15:0] _T_4480; // @[Mux.scala 31:69:@2146.4]
  wire  _T_4481; // @[OneHot.scala 66:30:@2147.4]
  wire  _T_4482; // @[OneHot.scala 66:30:@2148.4]
  wire  _T_4483; // @[OneHot.scala 66:30:@2149.4]
  wire  _T_4484; // @[OneHot.scala 66:30:@2150.4]
  wire  _T_4485; // @[OneHot.scala 66:30:@2151.4]
  wire  _T_4486; // @[OneHot.scala 66:30:@2152.4]
  wire  _T_4487; // @[OneHot.scala 66:30:@2153.4]
  wire  _T_4488; // @[OneHot.scala 66:30:@2154.4]
  wire  _T_4489; // @[OneHot.scala 66:30:@2155.4]
  wire  _T_4490; // @[OneHot.scala 66:30:@2156.4]
  wire  _T_4491; // @[OneHot.scala 66:30:@2157.4]
  wire  _T_4492; // @[OneHot.scala 66:30:@2158.4]
  wire  _T_4493; // @[OneHot.scala 66:30:@2159.4]
  wire  _T_4494; // @[OneHot.scala 66:30:@2160.4]
  wire  _T_4495; // @[OneHot.scala 66:30:@2161.4]
  wire  _T_4496; // @[OneHot.scala 66:30:@2162.4]
  wire [15:0] _T_4537; // @[Mux.scala 31:69:@2180.4]
  wire [15:0] _T_4538; // @[Mux.scala 31:69:@2181.4]
  wire [15:0] _T_4539; // @[Mux.scala 31:69:@2182.4]
  wire [15:0] _T_4540; // @[Mux.scala 31:69:@2183.4]
  wire [15:0] _T_4541; // @[Mux.scala 31:69:@2184.4]
  wire [15:0] _T_4542; // @[Mux.scala 31:69:@2185.4]
  wire [15:0] _T_4543; // @[Mux.scala 31:69:@2186.4]
  wire [15:0] _T_4544; // @[Mux.scala 31:69:@2187.4]
  wire [15:0] _T_4545; // @[Mux.scala 31:69:@2188.4]
  wire [15:0] _T_4546; // @[Mux.scala 31:69:@2189.4]
  wire [15:0] _T_4547; // @[Mux.scala 31:69:@2190.4]
  wire [15:0] _T_4548; // @[Mux.scala 31:69:@2191.4]
  wire [15:0] _T_4549; // @[Mux.scala 31:69:@2192.4]
  wire [15:0] _T_4550; // @[Mux.scala 31:69:@2193.4]
  wire [15:0] _T_4551; // @[Mux.scala 31:69:@2194.4]
  wire [15:0] _T_4552; // @[Mux.scala 31:69:@2195.4]
  wire  _T_4553; // @[OneHot.scala 66:30:@2196.4]
  wire  _T_4554; // @[OneHot.scala 66:30:@2197.4]
  wire  _T_4555; // @[OneHot.scala 66:30:@2198.4]
  wire  _T_4556; // @[OneHot.scala 66:30:@2199.4]
  wire  _T_4557; // @[OneHot.scala 66:30:@2200.4]
  wire  _T_4558; // @[OneHot.scala 66:30:@2201.4]
  wire  _T_4559; // @[OneHot.scala 66:30:@2202.4]
  wire  _T_4560; // @[OneHot.scala 66:30:@2203.4]
  wire  _T_4561; // @[OneHot.scala 66:30:@2204.4]
  wire  _T_4562; // @[OneHot.scala 66:30:@2205.4]
  wire  _T_4563; // @[OneHot.scala 66:30:@2206.4]
  wire  _T_4564; // @[OneHot.scala 66:30:@2207.4]
  wire  _T_4565; // @[OneHot.scala 66:30:@2208.4]
  wire  _T_4566; // @[OneHot.scala 66:30:@2209.4]
  wire  _T_4567; // @[OneHot.scala 66:30:@2210.4]
  wire  _T_4568; // @[OneHot.scala 66:30:@2211.4]
  wire [15:0] _T_4609; // @[Mux.scala 31:69:@2229.4]
  wire [15:0] _T_4610; // @[Mux.scala 31:69:@2230.4]
  wire [15:0] _T_4611; // @[Mux.scala 31:69:@2231.4]
  wire [15:0] _T_4612; // @[Mux.scala 31:69:@2232.4]
  wire [15:0] _T_4613; // @[Mux.scala 31:69:@2233.4]
  wire [15:0] _T_4614; // @[Mux.scala 31:69:@2234.4]
  wire [15:0] _T_4615; // @[Mux.scala 31:69:@2235.4]
  wire [15:0] _T_4616; // @[Mux.scala 31:69:@2236.4]
  wire [15:0] _T_4617; // @[Mux.scala 31:69:@2237.4]
  wire [15:0] _T_4618; // @[Mux.scala 31:69:@2238.4]
  wire [15:0] _T_4619; // @[Mux.scala 31:69:@2239.4]
  wire [15:0] _T_4620; // @[Mux.scala 31:69:@2240.4]
  wire [15:0] _T_4621; // @[Mux.scala 31:69:@2241.4]
  wire [15:0] _T_4622; // @[Mux.scala 31:69:@2242.4]
  wire [15:0] _T_4623; // @[Mux.scala 31:69:@2243.4]
  wire [15:0] _T_4624; // @[Mux.scala 31:69:@2244.4]
  wire  _T_4625; // @[OneHot.scala 66:30:@2245.4]
  wire  _T_4626; // @[OneHot.scala 66:30:@2246.4]
  wire  _T_4627; // @[OneHot.scala 66:30:@2247.4]
  wire  _T_4628; // @[OneHot.scala 66:30:@2248.4]
  wire  _T_4629; // @[OneHot.scala 66:30:@2249.4]
  wire  _T_4630; // @[OneHot.scala 66:30:@2250.4]
  wire  _T_4631; // @[OneHot.scala 66:30:@2251.4]
  wire  _T_4632; // @[OneHot.scala 66:30:@2252.4]
  wire  _T_4633; // @[OneHot.scala 66:30:@2253.4]
  wire  _T_4634; // @[OneHot.scala 66:30:@2254.4]
  wire  _T_4635; // @[OneHot.scala 66:30:@2255.4]
  wire  _T_4636; // @[OneHot.scala 66:30:@2256.4]
  wire  _T_4637; // @[OneHot.scala 66:30:@2257.4]
  wire  _T_4638; // @[OneHot.scala 66:30:@2258.4]
  wire  _T_4639; // @[OneHot.scala 66:30:@2259.4]
  wire  _T_4640; // @[OneHot.scala 66:30:@2260.4]
  wire [15:0] _T_4681; // @[Mux.scala 31:69:@2278.4]
  wire [15:0] _T_4682; // @[Mux.scala 31:69:@2279.4]
  wire [15:0] _T_4683; // @[Mux.scala 31:69:@2280.4]
  wire [15:0] _T_4684; // @[Mux.scala 31:69:@2281.4]
  wire [15:0] _T_4685; // @[Mux.scala 31:69:@2282.4]
  wire [15:0] _T_4686; // @[Mux.scala 31:69:@2283.4]
  wire [15:0] _T_4687; // @[Mux.scala 31:69:@2284.4]
  wire [15:0] _T_4688; // @[Mux.scala 31:69:@2285.4]
  wire [15:0] _T_4689; // @[Mux.scala 31:69:@2286.4]
  wire [15:0] _T_4690; // @[Mux.scala 31:69:@2287.4]
  wire [15:0] _T_4691; // @[Mux.scala 31:69:@2288.4]
  wire [15:0] _T_4692; // @[Mux.scala 31:69:@2289.4]
  wire [15:0] _T_4693; // @[Mux.scala 31:69:@2290.4]
  wire [15:0] _T_4694; // @[Mux.scala 31:69:@2291.4]
  wire [15:0] _T_4695; // @[Mux.scala 31:69:@2292.4]
  wire [15:0] _T_4696; // @[Mux.scala 31:69:@2293.4]
  wire  _T_4697; // @[OneHot.scala 66:30:@2294.4]
  wire  _T_4698; // @[OneHot.scala 66:30:@2295.4]
  wire  _T_4699; // @[OneHot.scala 66:30:@2296.4]
  wire  _T_4700; // @[OneHot.scala 66:30:@2297.4]
  wire  _T_4701; // @[OneHot.scala 66:30:@2298.4]
  wire  _T_4702; // @[OneHot.scala 66:30:@2299.4]
  wire  _T_4703; // @[OneHot.scala 66:30:@2300.4]
  wire  _T_4704; // @[OneHot.scala 66:30:@2301.4]
  wire  _T_4705; // @[OneHot.scala 66:30:@2302.4]
  wire  _T_4706; // @[OneHot.scala 66:30:@2303.4]
  wire  _T_4707; // @[OneHot.scala 66:30:@2304.4]
  wire  _T_4708; // @[OneHot.scala 66:30:@2305.4]
  wire  _T_4709; // @[OneHot.scala 66:30:@2306.4]
  wire  _T_4710; // @[OneHot.scala 66:30:@2307.4]
  wire  _T_4711; // @[OneHot.scala 66:30:@2308.4]
  wire  _T_4712; // @[OneHot.scala 66:30:@2309.4]
  wire [15:0] _T_4753; // @[Mux.scala 31:69:@2327.4]
  wire [15:0] _T_4754; // @[Mux.scala 31:69:@2328.4]
  wire [15:0] _T_4755; // @[Mux.scala 31:69:@2329.4]
  wire [15:0] _T_4756; // @[Mux.scala 31:69:@2330.4]
  wire [15:0] _T_4757; // @[Mux.scala 31:69:@2331.4]
  wire [15:0] _T_4758; // @[Mux.scala 31:69:@2332.4]
  wire [15:0] _T_4759; // @[Mux.scala 31:69:@2333.4]
  wire [15:0] _T_4760; // @[Mux.scala 31:69:@2334.4]
  wire [15:0] _T_4761; // @[Mux.scala 31:69:@2335.4]
  wire [15:0] _T_4762; // @[Mux.scala 31:69:@2336.4]
  wire [15:0] _T_4763; // @[Mux.scala 31:69:@2337.4]
  wire [15:0] _T_4764; // @[Mux.scala 31:69:@2338.4]
  wire [15:0] _T_4765; // @[Mux.scala 31:69:@2339.4]
  wire [15:0] _T_4766; // @[Mux.scala 31:69:@2340.4]
  wire [15:0] _T_4767; // @[Mux.scala 31:69:@2341.4]
  wire [15:0] _T_4768; // @[Mux.scala 31:69:@2342.4]
  wire  _T_4769; // @[OneHot.scala 66:30:@2343.4]
  wire  _T_4770; // @[OneHot.scala 66:30:@2344.4]
  wire  _T_4771; // @[OneHot.scala 66:30:@2345.4]
  wire  _T_4772; // @[OneHot.scala 66:30:@2346.4]
  wire  _T_4773; // @[OneHot.scala 66:30:@2347.4]
  wire  _T_4774; // @[OneHot.scala 66:30:@2348.4]
  wire  _T_4775; // @[OneHot.scala 66:30:@2349.4]
  wire  _T_4776; // @[OneHot.scala 66:30:@2350.4]
  wire  _T_4777; // @[OneHot.scala 66:30:@2351.4]
  wire  _T_4778; // @[OneHot.scala 66:30:@2352.4]
  wire  _T_4779; // @[OneHot.scala 66:30:@2353.4]
  wire  _T_4780; // @[OneHot.scala 66:30:@2354.4]
  wire  _T_4781; // @[OneHot.scala 66:30:@2355.4]
  wire  _T_4782; // @[OneHot.scala 66:30:@2356.4]
  wire  _T_4783; // @[OneHot.scala 66:30:@2357.4]
  wire  _T_4784; // @[OneHot.scala 66:30:@2358.4]
  wire [15:0] _T_4825; // @[Mux.scala 31:69:@2376.4]
  wire [15:0] _T_4826; // @[Mux.scala 31:69:@2377.4]
  wire [15:0] _T_4827; // @[Mux.scala 31:69:@2378.4]
  wire [15:0] _T_4828; // @[Mux.scala 31:69:@2379.4]
  wire [15:0] _T_4829; // @[Mux.scala 31:69:@2380.4]
  wire [15:0] _T_4830; // @[Mux.scala 31:69:@2381.4]
  wire [15:0] _T_4831; // @[Mux.scala 31:69:@2382.4]
  wire [15:0] _T_4832; // @[Mux.scala 31:69:@2383.4]
  wire [15:0] _T_4833; // @[Mux.scala 31:69:@2384.4]
  wire [15:0] _T_4834; // @[Mux.scala 31:69:@2385.4]
  wire [15:0] _T_4835; // @[Mux.scala 31:69:@2386.4]
  wire [15:0] _T_4836; // @[Mux.scala 31:69:@2387.4]
  wire [15:0] _T_4837; // @[Mux.scala 31:69:@2388.4]
  wire [15:0] _T_4838; // @[Mux.scala 31:69:@2389.4]
  wire [15:0] _T_4839; // @[Mux.scala 31:69:@2390.4]
  wire [15:0] _T_4840; // @[Mux.scala 31:69:@2391.4]
  wire  _T_4841; // @[OneHot.scala 66:30:@2392.4]
  wire  _T_4842; // @[OneHot.scala 66:30:@2393.4]
  wire  _T_4843; // @[OneHot.scala 66:30:@2394.4]
  wire  _T_4844; // @[OneHot.scala 66:30:@2395.4]
  wire  _T_4845; // @[OneHot.scala 66:30:@2396.4]
  wire  _T_4846; // @[OneHot.scala 66:30:@2397.4]
  wire  _T_4847; // @[OneHot.scala 66:30:@2398.4]
  wire  _T_4848; // @[OneHot.scala 66:30:@2399.4]
  wire  _T_4849; // @[OneHot.scala 66:30:@2400.4]
  wire  _T_4850; // @[OneHot.scala 66:30:@2401.4]
  wire  _T_4851; // @[OneHot.scala 66:30:@2402.4]
  wire  _T_4852; // @[OneHot.scala 66:30:@2403.4]
  wire  _T_4853; // @[OneHot.scala 66:30:@2404.4]
  wire  _T_4854; // @[OneHot.scala 66:30:@2405.4]
  wire  _T_4855; // @[OneHot.scala 66:30:@2406.4]
  wire  _T_4856; // @[OneHot.scala 66:30:@2407.4]
  wire [15:0] _T_4897; // @[Mux.scala 31:69:@2425.4]
  wire [15:0] _T_4898; // @[Mux.scala 31:69:@2426.4]
  wire [15:0] _T_4899; // @[Mux.scala 31:69:@2427.4]
  wire [15:0] _T_4900; // @[Mux.scala 31:69:@2428.4]
  wire [15:0] _T_4901; // @[Mux.scala 31:69:@2429.4]
  wire [15:0] _T_4902; // @[Mux.scala 31:69:@2430.4]
  wire [15:0] _T_4903; // @[Mux.scala 31:69:@2431.4]
  wire [15:0] _T_4904; // @[Mux.scala 31:69:@2432.4]
  wire [15:0] _T_4905; // @[Mux.scala 31:69:@2433.4]
  wire [15:0] _T_4906; // @[Mux.scala 31:69:@2434.4]
  wire [15:0] _T_4907; // @[Mux.scala 31:69:@2435.4]
  wire [15:0] _T_4908; // @[Mux.scala 31:69:@2436.4]
  wire [15:0] _T_4909; // @[Mux.scala 31:69:@2437.4]
  wire [15:0] _T_4910; // @[Mux.scala 31:69:@2438.4]
  wire [15:0] _T_4911; // @[Mux.scala 31:69:@2439.4]
  wire [15:0] _T_4912; // @[Mux.scala 31:69:@2440.4]
  wire  _T_4913; // @[OneHot.scala 66:30:@2441.4]
  wire  _T_4914; // @[OneHot.scala 66:30:@2442.4]
  wire  _T_4915; // @[OneHot.scala 66:30:@2443.4]
  wire  _T_4916; // @[OneHot.scala 66:30:@2444.4]
  wire  _T_4917; // @[OneHot.scala 66:30:@2445.4]
  wire  _T_4918; // @[OneHot.scala 66:30:@2446.4]
  wire  _T_4919; // @[OneHot.scala 66:30:@2447.4]
  wire  _T_4920; // @[OneHot.scala 66:30:@2448.4]
  wire  _T_4921; // @[OneHot.scala 66:30:@2449.4]
  wire  _T_4922; // @[OneHot.scala 66:30:@2450.4]
  wire  _T_4923; // @[OneHot.scala 66:30:@2451.4]
  wire  _T_4924; // @[OneHot.scala 66:30:@2452.4]
  wire  _T_4925; // @[OneHot.scala 66:30:@2453.4]
  wire  _T_4926; // @[OneHot.scala 66:30:@2454.4]
  wire  _T_4927; // @[OneHot.scala 66:30:@2455.4]
  wire  _T_4928; // @[OneHot.scala 66:30:@2456.4]
  wire [15:0] _T_4969; // @[Mux.scala 31:69:@2474.4]
  wire [15:0] _T_4970; // @[Mux.scala 31:69:@2475.4]
  wire [15:0] _T_4971; // @[Mux.scala 31:69:@2476.4]
  wire [15:0] _T_4972; // @[Mux.scala 31:69:@2477.4]
  wire [15:0] _T_4973; // @[Mux.scala 31:69:@2478.4]
  wire [15:0] _T_4974; // @[Mux.scala 31:69:@2479.4]
  wire [15:0] _T_4975; // @[Mux.scala 31:69:@2480.4]
  wire [15:0] _T_4976; // @[Mux.scala 31:69:@2481.4]
  wire [15:0] _T_4977; // @[Mux.scala 31:69:@2482.4]
  wire [15:0] _T_4978; // @[Mux.scala 31:69:@2483.4]
  wire [15:0] _T_4979; // @[Mux.scala 31:69:@2484.4]
  wire [15:0] _T_4980; // @[Mux.scala 31:69:@2485.4]
  wire [15:0] _T_4981; // @[Mux.scala 31:69:@2486.4]
  wire [15:0] _T_4982; // @[Mux.scala 31:69:@2487.4]
  wire [15:0] _T_4983; // @[Mux.scala 31:69:@2488.4]
  wire [15:0] _T_4984; // @[Mux.scala 31:69:@2489.4]
  wire  _T_4985; // @[OneHot.scala 66:30:@2490.4]
  wire  _T_4986; // @[OneHot.scala 66:30:@2491.4]
  wire  _T_4987; // @[OneHot.scala 66:30:@2492.4]
  wire  _T_4988; // @[OneHot.scala 66:30:@2493.4]
  wire  _T_4989; // @[OneHot.scala 66:30:@2494.4]
  wire  _T_4990; // @[OneHot.scala 66:30:@2495.4]
  wire  _T_4991; // @[OneHot.scala 66:30:@2496.4]
  wire  _T_4992; // @[OneHot.scala 66:30:@2497.4]
  wire  _T_4993; // @[OneHot.scala 66:30:@2498.4]
  wire  _T_4994; // @[OneHot.scala 66:30:@2499.4]
  wire  _T_4995; // @[OneHot.scala 66:30:@2500.4]
  wire  _T_4996; // @[OneHot.scala 66:30:@2501.4]
  wire  _T_4997; // @[OneHot.scala 66:30:@2502.4]
  wire  _T_4998; // @[OneHot.scala 66:30:@2503.4]
  wire  _T_4999; // @[OneHot.scala 66:30:@2504.4]
  wire  _T_5000; // @[OneHot.scala 66:30:@2505.4]
  wire [15:0] _T_5041; // @[Mux.scala 31:69:@2523.4]
  wire [15:0] _T_5042; // @[Mux.scala 31:69:@2524.4]
  wire [15:0] _T_5043; // @[Mux.scala 31:69:@2525.4]
  wire [15:0] _T_5044; // @[Mux.scala 31:69:@2526.4]
  wire [15:0] _T_5045; // @[Mux.scala 31:69:@2527.4]
  wire [15:0] _T_5046; // @[Mux.scala 31:69:@2528.4]
  wire [15:0] _T_5047; // @[Mux.scala 31:69:@2529.4]
  wire [15:0] _T_5048; // @[Mux.scala 31:69:@2530.4]
  wire [15:0] _T_5049; // @[Mux.scala 31:69:@2531.4]
  wire [15:0] _T_5050; // @[Mux.scala 31:69:@2532.4]
  wire [15:0] _T_5051; // @[Mux.scala 31:69:@2533.4]
  wire [15:0] _T_5052; // @[Mux.scala 31:69:@2534.4]
  wire [15:0] _T_5053; // @[Mux.scala 31:69:@2535.4]
  wire [15:0] _T_5054; // @[Mux.scala 31:69:@2536.4]
  wire [15:0] _T_5055; // @[Mux.scala 31:69:@2537.4]
  wire [15:0] _T_5056; // @[Mux.scala 31:69:@2538.4]
  wire  _T_5057; // @[OneHot.scala 66:30:@2539.4]
  wire  _T_5058; // @[OneHot.scala 66:30:@2540.4]
  wire  _T_5059; // @[OneHot.scala 66:30:@2541.4]
  wire  _T_5060; // @[OneHot.scala 66:30:@2542.4]
  wire  _T_5061; // @[OneHot.scala 66:30:@2543.4]
  wire  _T_5062; // @[OneHot.scala 66:30:@2544.4]
  wire  _T_5063; // @[OneHot.scala 66:30:@2545.4]
  wire  _T_5064; // @[OneHot.scala 66:30:@2546.4]
  wire  _T_5065; // @[OneHot.scala 66:30:@2547.4]
  wire  _T_5066; // @[OneHot.scala 66:30:@2548.4]
  wire  _T_5067; // @[OneHot.scala 66:30:@2549.4]
  wire  _T_5068; // @[OneHot.scala 66:30:@2550.4]
  wire  _T_5069; // @[OneHot.scala 66:30:@2551.4]
  wire  _T_5070; // @[OneHot.scala 66:30:@2552.4]
  wire  _T_5071; // @[OneHot.scala 66:30:@2553.4]
  wire  _T_5072; // @[OneHot.scala 66:30:@2554.4]
  wire [15:0] _T_5113; // @[Mux.scala 31:69:@2572.4]
  wire [15:0] _T_5114; // @[Mux.scala 31:69:@2573.4]
  wire [15:0] _T_5115; // @[Mux.scala 31:69:@2574.4]
  wire [15:0] _T_5116; // @[Mux.scala 31:69:@2575.4]
  wire [15:0] _T_5117; // @[Mux.scala 31:69:@2576.4]
  wire [15:0] _T_5118; // @[Mux.scala 31:69:@2577.4]
  wire [15:0] _T_5119; // @[Mux.scala 31:69:@2578.4]
  wire [15:0] _T_5120; // @[Mux.scala 31:69:@2579.4]
  wire [15:0] _T_5121; // @[Mux.scala 31:69:@2580.4]
  wire [15:0] _T_5122; // @[Mux.scala 31:69:@2581.4]
  wire [15:0] _T_5123; // @[Mux.scala 31:69:@2582.4]
  wire [15:0] _T_5124; // @[Mux.scala 31:69:@2583.4]
  wire [15:0] _T_5125; // @[Mux.scala 31:69:@2584.4]
  wire [15:0] _T_5126; // @[Mux.scala 31:69:@2585.4]
  wire [15:0] _T_5127; // @[Mux.scala 31:69:@2586.4]
  wire [15:0] _T_5128; // @[Mux.scala 31:69:@2587.4]
  wire  _T_5129; // @[OneHot.scala 66:30:@2588.4]
  wire  _T_5130; // @[OneHot.scala 66:30:@2589.4]
  wire  _T_5131; // @[OneHot.scala 66:30:@2590.4]
  wire  _T_5132; // @[OneHot.scala 66:30:@2591.4]
  wire  _T_5133; // @[OneHot.scala 66:30:@2592.4]
  wire  _T_5134; // @[OneHot.scala 66:30:@2593.4]
  wire  _T_5135; // @[OneHot.scala 66:30:@2594.4]
  wire  _T_5136; // @[OneHot.scala 66:30:@2595.4]
  wire  _T_5137; // @[OneHot.scala 66:30:@2596.4]
  wire  _T_5138; // @[OneHot.scala 66:30:@2597.4]
  wire  _T_5139; // @[OneHot.scala 66:30:@2598.4]
  wire  _T_5140; // @[OneHot.scala 66:30:@2599.4]
  wire  _T_5141; // @[OneHot.scala 66:30:@2600.4]
  wire  _T_5142; // @[OneHot.scala 66:30:@2601.4]
  wire  _T_5143; // @[OneHot.scala 66:30:@2602.4]
  wire  _T_5144; // @[OneHot.scala 66:30:@2603.4]
  wire [15:0] _T_5185; // @[Mux.scala 31:69:@2621.4]
  wire [15:0] _T_5186; // @[Mux.scala 31:69:@2622.4]
  wire [15:0] _T_5187; // @[Mux.scala 31:69:@2623.4]
  wire [15:0] _T_5188; // @[Mux.scala 31:69:@2624.4]
  wire [15:0] _T_5189; // @[Mux.scala 31:69:@2625.4]
  wire [15:0] _T_5190; // @[Mux.scala 31:69:@2626.4]
  wire [15:0] _T_5191; // @[Mux.scala 31:69:@2627.4]
  wire [15:0] _T_5192; // @[Mux.scala 31:69:@2628.4]
  wire [15:0] _T_5193; // @[Mux.scala 31:69:@2629.4]
  wire [15:0] _T_5194; // @[Mux.scala 31:69:@2630.4]
  wire [15:0] _T_5195; // @[Mux.scala 31:69:@2631.4]
  wire [15:0] _T_5196; // @[Mux.scala 31:69:@2632.4]
  wire [15:0] _T_5197; // @[Mux.scala 31:69:@2633.4]
  wire [15:0] _T_5198; // @[Mux.scala 31:69:@2634.4]
  wire [15:0] _T_5199; // @[Mux.scala 31:69:@2635.4]
  wire [15:0] _T_5200; // @[Mux.scala 31:69:@2636.4]
  wire  _T_5201; // @[OneHot.scala 66:30:@2637.4]
  wire  _T_5202; // @[OneHot.scala 66:30:@2638.4]
  wire  _T_5203; // @[OneHot.scala 66:30:@2639.4]
  wire  _T_5204; // @[OneHot.scala 66:30:@2640.4]
  wire  _T_5205; // @[OneHot.scala 66:30:@2641.4]
  wire  _T_5206; // @[OneHot.scala 66:30:@2642.4]
  wire  _T_5207; // @[OneHot.scala 66:30:@2643.4]
  wire  _T_5208; // @[OneHot.scala 66:30:@2644.4]
  wire  _T_5209; // @[OneHot.scala 66:30:@2645.4]
  wire  _T_5210; // @[OneHot.scala 66:30:@2646.4]
  wire  _T_5211; // @[OneHot.scala 66:30:@2647.4]
  wire  _T_5212; // @[OneHot.scala 66:30:@2648.4]
  wire  _T_5213; // @[OneHot.scala 66:30:@2649.4]
  wire  _T_5214; // @[OneHot.scala 66:30:@2650.4]
  wire  _T_5215; // @[OneHot.scala 66:30:@2651.4]
  wire  _T_5216; // @[OneHot.scala 66:30:@2652.4]
  wire [15:0] _T_5257; // @[Mux.scala 31:69:@2670.4]
  wire [15:0] _T_5258; // @[Mux.scala 31:69:@2671.4]
  wire [15:0] _T_5259; // @[Mux.scala 31:69:@2672.4]
  wire [15:0] _T_5260; // @[Mux.scala 31:69:@2673.4]
  wire [15:0] _T_5261; // @[Mux.scala 31:69:@2674.4]
  wire [15:0] _T_5262; // @[Mux.scala 31:69:@2675.4]
  wire [15:0] _T_5263; // @[Mux.scala 31:69:@2676.4]
  wire [15:0] _T_5264; // @[Mux.scala 31:69:@2677.4]
  wire [15:0] _T_5265; // @[Mux.scala 31:69:@2678.4]
  wire [15:0] _T_5266; // @[Mux.scala 31:69:@2679.4]
  wire [15:0] _T_5267; // @[Mux.scala 31:69:@2680.4]
  wire [15:0] _T_5268; // @[Mux.scala 31:69:@2681.4]
  wire [15:0] _T_5269; // @[Mux.scala 31:69:@2682.4]
  wire [15:0] _T_5270; // @[Mux.scala 31:69:@2683.4]
  wire [15:0] _T_5271; // @[Mux.scala 31:69:@2684.4]
  wire [15:0] _T_5272; // @[Mux.scala 31:69:@2685.4]
  wire  _T_5273; // @[OneHot.scala 66:30:@2686.4]
  wire  _T_5274; // @[OneHot.scala 66:30:@2687.4]
  wire  _T_5275; // @[OneHot.scala 66:30:@2688.4]
  wire  _T_5276; // @[OneHot.scala 66:30:@2689.4]
  wire  _T_5277; // @[OneHot.scala 66:30:@2690.4]
  wire  _T_5278; // @[OneHot.scala 66:30:@2691.4]
  wire  _T_5279; // @[OneHot.scala 66:30:@2692.4]
  wire  _T_5280; // @[OneHot.scala 66:30:@2693.4]
  wire  _T_5281; // @[OneHot.scala 66:30:@2694.4]
  wire  _T_5282; // @[OneHot.scala 66:30:@2695.4]
  wire  _T_5283; // @[OneHot.scala 66:30:@2696.4]
  wire  _T_5284; // @[OneHot.scala 66:30:@2697.4]
  wire  _T_5285; // @[OneHot.scala 66:30:@2698.4]
  wire  _T_5286; // @[OneHot.scala 66:30:@2699.4]
  wire  _T_5287; // @[OneHot.scala 66:30:@2700.4]
  wire  _T_5288; // @[OneHot.scala 66:30:@2701.4]
  wire [15:0] _T_5329; // @[Mux.scala 31:69:@2719.4]
  wire [15:0] _T_5330; // @[Mux.scala 31:69:@2720.4]
  wire [15:0] _T_5331; // @[Mux.scala 31:69:@2721.4]
  wire [15:0] _T_5332; // @[Mux.scala 31:69:@2722.4]
  wire [15:0] _T_5333; // @[Mux.scala 31:69:@2723.4]
  wire [15:0] _T_5334; // @[Mux.scala 31:69:@2724.4]
  wire [15:0] _T_5335; // @[Mux.scala 31:69:@2725.4]
  wire [15:0] _T_5336; // @[Mux.scala 31:69:@2726.4]
  wire [15:0] _T_5337; // @[Mux.scala 31:69:@2727.4]
  wire [15:0] _T_5338; // @[Mux.scala 31:69:@2728.4]
  wire [15:0] _T_5339; // @[Mux.scala 31:69:@2729.4]
  wire [15:0] _T_5340; // @[Mux.scala 31:69:@2730.4]
  wire [15:0] _T_5341; // @[Mux.scala 31:69:@2731.4]
  wire [15:0] _T_5342; // @[Mux.scala 31:69:@2732.4]
  wire [15:0] _T_5343; // @[Mux.scala 31:69:@2733.4]
  wire [15:0] _T_5344; // @[Mux.scala 31:69:@2734.4]
  wire  _T_5345; // @[OneHot.scala 66:30:@2735.4]
  wire  _T_5346; // @[OneHot.scala 66:30:@2736.4]
  wire  _T_5347; // @[OneHot.scala 66:30:@2737.4]
  wire  _T_5348; // @[OneHot.scala 66:30:@2738.4]
  wire  _T_5349; // @[OneHot.scala 66:30:@2739.4]
  wire  _T_5350; // @[OneHot.scala 66:30:@2740.4]
  wire  _T_5351; // @[OneHot.scala 66:30:@2741.4]
  wire  _T_5352; // @[OneHot.scala 66:30:@2742.4]
  wire  _T_5353; // @[OneHot.scala 66:30:@2743.4]
  wire  _T_5354; // @[OneHot.scala 66:30:@2744.4]
  wire  _T_5355; // @[OneHot.scala 66:30:@2745.4]
  wire  _T_5356; // @[OneHot.scala 66:30:@2746.4]
  wire  _T_5357; // @[OneHot.scala 66:30:@2747.4]
  wire  _T_5358; // @[OneHot.scala 66:30:@2748.4]
  wire  _T_5359; // @[OneHot.scala 66:30:@2749.4]
  wire  _T_5360; // @[OneHot.scala 66:30:@2750.4]
  wire [15:0] _T_5401; // @[Mux.scala 31:69:@2768.4]
  wire [15:0] _T_5402; // @[Mux.scala 31:69:@2769.4]
  wire [15:0] _T_5403; // @[Mux.scala 31:69:@2770.4]
  wire [15:0] _T_5404; // @[Mux.scala 31:69:@2771.4]
  wire [15:0] _T_5405; // @[Mux.scala 31:69:@2772.4]
  wire [15:0] _T_5406; // @[Mux.scala 31:69:@2773.4]
  wire [15:0] _T_5407; // @[Mux.scala 31:69:@2774.4]
  wire [15:0] _T_5408; // @[Mux.scala 31:69:@2775.4]
  wire [15:0] _T_5409; // @[Mux.scala 31:69:@2776.4]
  wire [15:0] _T_5410; // @[Mux.scala 31:69:@2777.4]
  wire [15:0] _T_5411; // @[Mux.scala 31:69:@2778.4]
  wire [15:0] _T_5412; // @[Mux.scala 31:69:@2779.4]
  wire [15:0] _T_5413; // @[Mux.scala 31:69:@2780.4]
  wire [15:0] _T_5414; // @[Mux.scala 31:69:@2781.4]
  wire [15:0] _T_5415; // @[Mux.scala 31:69:@2782.4]
  wire [15:0] _T_5416; // @[Mux.scala 31:69:@2783.4]
  wire  _T_5417; // @[OneHot.scala 66:30:@2784.4]
  wire  _T_5418; // @[OneHot.scala 66:30:@2785.4]
  wire  _T_5419; // @[OneHot.scala 66:30:@2786.4]
  wire  _T_5420; // @[OneHot.scala 66:30:@2787.4]
  wire  _T_5421; // @[OneHot.scala 66:30:@2788.4]
  wire  _T_5422; // @[OneHot.scala 66:30:@2789.4]
  wire  _T_5423; // @[OneHot.scala 66:30:@2790.4]
  wire  _T_5424; // @[OneHot.scala 66:30:@2791.4]
  wire  _T_5425; // @[OneHot.scala 66:30:@2792.4]
  wire  _T_5426; // @[OneHot.scala 66:30:@2793.4]
  wire  _T_5427; // @[OneHot.scala 66:30:@2794.4]
  wire  _T_5428; // @[OneHot.scala 66:30:@2795.4]
  wire  _T_5429; // @[OneHot.scala 66:30:@2796.4]
  wire  _T_5430; // @[OneHot.scala 66:30:@2797.4]
  wire  _T_5431; // @[OneHot.scala 66:30:@2798.4]
  wire  _T_5432; // @[OneHot.scala 66:30:@2799.4]
  wire [7:0] _T_5497; // @[Mux.scala 19:72:@2823.4]
  wire [15:0] _T_5505; // @[Mux.scala 19:72:@2831.4]
  wire [15:0] _T_5507; // @[Mux.scala 19:72:@2832.4]
  wire [7:0] _T_5514; // @[Mux.scala 19:72:@2839.4]
  wire [15:0] _T_5522; // @[Mux.scala 19:72:@2847.4]
  wire [15:0] _T_5524; // @[Mux.scala 19:72:@2848.4]
  wire [7:0] _T_5531; // @[Mux.scala 19:72:@2855.4]
  wire [15:0] _T_5539; // @[Mux.scala 19:72:@2863.4]
  wire [15:0] _T_5541; // @[Mux.scala 19:72:@2864.4]
  wire [7:0] _T_5548; // @[Mux.scala 19:72:@2871.4]
  wire [15:0] _T_5556; // @[Mux.scala 19:72:@2879.4]
  wire [15:0] _T_5558; // @[Mux.scala 19:72:@2880.4]
  wire [7:0] _T_5565; // @[Mux.scala 19:72:@2887.4]
  wire [15:0] _T_5573; // @[Mux.scala 19:72:@2895.4]
  wire [15:0] _T_5575; // @[Mux.scala 19:72:@2896.4]
  wire [7:0] _T_5582; // @[Mux.scala 19:72:@2903.4]
  wire [15:0] _T_5590; // @[Mux.scala 19:72:@2911.4]
  wire [15:0] _T_5592; // @[Mux.scala 19:72:@2912.4]
  wire [7:0] _T_5599; // @[Mux.scala 19:72:@2919.4]
  wire [15:0] _T_5607; // @[Mux.scala 19:72:@2927.4]
  wire [15:0] _T_5609; // @[Mux.scala 19:72:@2928.4]
  wire [7:0] _T_5616; // @[Mux.scala 19:72:@2935.4]
  wire [15:0] _T_5624; // @[Mux.scala 19:72:@2943.4]
  wire [15:0] _T_5626; // @[Mux.scala 19:72:@2944.4]
  wire [7:0] _T_5633; // @[Mux.scala 19:72:@2951.4]
  wire [15:0] _T_5641; // @[Mux.scala 19:72:@2959.4]
  wire [15:0] _T_5643; // @[Mux.scala 19:72:@2960.4]
  wire [7:0] _T_5650; // @[Mux.scala 19:72:@2967.4]
  wire [15:0] _T_5658; // @[Mux.scala 19:72:@2975.4]
  wire [15:0] _T_5660; // @[Mux.scala 19:72:@2976.4]
  wire [7:0] _T_5667; // @[Mux.scala 19:72:@2983.4]
  wire [15:0] _T_5675; // @[Mux.scala 19:72:@2991.4]
  wire [15:0] _T_5677; // @[Mux.scala 19:72:@2992.4]
  wire [7:0] _T_5684; // @[Mux.scala 19:72:@2999.4]
  wire [15:0] _T_5692; // @[Mux.scala 19:72:@3007.4]
  wire [15:0] _T_5694; // @[Mux.scala 19:72:@3008.4]
  wire [7:0] _T_5701; // @[Mux.scala 19:72:@3015.4]
  wire [15:0] _T_5709; // @[Mux.scala 19:72:@3023.4]
  wire [15:0] _T_5711; // @[Mux.scala 19:72:@3024.4]
  wire [7:0] _T_5718; // @[Mux.scala 19:72:@3031.4]
  wire [15:0] _T_5726; // @[Mux.scala 19:72:@3039.4]
  wire [15:0] _T_5728; // @[Mux.scala 19:72:@3040.4]
  wire [7:0] _T_5735; // @[Mux.scala 19:72:@3047.4]
  wire [15:0] _T_5743; // @[Mux.scala 19:72:@3055.4]
  wire [15:0] _T_5745; // @[Mux.scala 19:72:@3056.4]
  wire [7:0] _T_5752; // @[Mux.scala 19:72:@3063.4]
  wire [15:0] _T_5760; // @[Mux.scala 19:72:@3071.4]
  wire [15:0] _T_5762; // @[Mux.scala 19:72:@3072.4]
  wire [15:0] _T_5763; // @[Mux.scala 19:72:@3073.4]
  wire [15:0] _T_5764; // @[Mux.scala 19:72:@3074.4]
  wire [15:0] _T_5765; // @[Mux.scala 19:72:@3075.4]
  wire [15:0] _T_5766; // @[Mux.scala 19:72:@3076.4]
  wire [15:0] _T_5767; // @[Mux.scala 19:72:@3077.4]
  wire [15:0] _T_5768; // @[Mux.scala 19:72:@3078.4]
  wire [15:0] _T_5769; // @[Mux.scala 19:72:@3079.4]
  wire [15:0] _T_5770; // @[Mux.scala 19:72:@3080.4]
  wire [15:0] _T_5771; // @[Mux.scala 19:72:@3081.4]
  wire [15:0] _T_5772; // @[Mux.scala 19:72:@3082.4]
  wire [15:0] _T_5773; // @[Mux.scala 19:72:@3083.4]
  wire [15:0] _T_5774; // @[Mux.scala 19:72:@3084.4]
  wire [15:0] _T_5775; // @[Mux.scala 19:72:@3085.4]
  wire [15:0] _T_5776; // @[Mux.scala 19:72:@3086.4]
  wire [15:0] _T_5777; // @[Mux.scala 19:72:@3087.4]
  wire  inputAddrPriorityPorts_0_0; // @[Mux.scala 19:72:@3091.4]
  wire  inputAddrPriorityPorts_0_1; // @[Mux.scala 19:72:@3093.4]
  wire  inputAddrPriorityPorts_0_2; // @[Mux.scala 19:72:@3095.4]
  wire  inputAddrPriorityPorts_0_3; // @[Mux.scala 19:72:@3097.4]
  wire  inputAddrPriorityPorts_0_4; // @[Mux.scala 19:72:@3099.4]
  wire  inputAddrPriorityPorts_0_5; // @[Mux.scala 19:72:@3101.4]
  wire  inputAddrPriorityPorts_0_6; // @[Mux.scala 19:72:@3103.4]
  wire  inputAddrPriorityPorts_0_7; // @[Mux.scala 19:72:@3105.4]
  wire  inputAddrPriorityPorts_0_8; // @[Mux.scala 19:72:@3107.4]
  wire  inputAddrPriorityPorts_0_9; // @[Mux.scala 19:72:@3109.4]
  wire  inputAddrPriorityPorts_0_10; // @[Mux.scala 19:72:@3111.4]
  wire  inputAddrPriorityPorts_0_11; // @[Mux.scala 19:72:@3113.4]
  wire  inputAddrPriorityPorts_0_12; // @[Mux.scala 19:72:@3115.4]
  wire  inputAddrPriorityPorts_0_13; // @[Mux.scala 19:72:@3117.4]
  wire  inputAddrPriorityPorts_0_14; // @[Mux.scala 19:72:@3119.4]
  wire  inputAddrPriorityPorts_0_15; // @[Mux.scala 19:72:@3121.4]
  wire [15:0] _T_5979; // @[Mux.scala 31:69:@3175.4]
  wire [15:0] _T_5980; // @[Mux.scala 31:69:@3176.4]
  wire [15:0] _T_5981; // @[Mux.scala 31:69:@3177.4]
  wire [15:0] _T_5982; // @[Mux.scala 31:69:@3178.4]
  wire [15:0] _T_5983; // @[Mux.scala 31:69:@3179.4]
  wire [15:0] _T_5984; // @[Mux.scala 31:69:@3180.4]
  wire [15:0] _T_5985; // @[Mux.scala 31:69:@3181.4]
  wire [15:0] _T_5986; // @[Mux.scala 31:69:@3182.4]
  wire [15:0] _T_5987; // @[Mux.scala 31:69:@3183.4]
  wire [15:0] _T_5988; // @[Mux.scala 31:69:@3184.4]
  wire [15:0] _T_5989; // @[Mux.scala 31:69:@3185.4]
  wire [15:0] _T_5990; // @[Mux.scala 31:69:@3186.4]
  wire [15:0] _T_5991; // @[Mux.scala 31:69:@3187.4]
  wire [15:0] _T_5992; // @[Mux.scala 31:69:@3188.4]
  wire [15:0] _T_5993; // @[Mux.scala 31:69:@3189.4]
  wire [15:0] _T_5994; // @[Mux.scala 31:69:@3190.4]
  wire  _T_5995; // @[OneHot.scala 66:30:@3191.4]
  wire  _T_5996; // @[OneHot.scala 66:30:@3192.4]
  wire  _T_5997; // @[OneHot.scala 66:30:@3193.4]
  wire  _T_5998; // @[OneHot.scala 66:30:@3194.4]
  wire  _T_5999; // @[OneHot.scala 66:30:@3195.4]
  wire  _T_6000; // @[OneHot.scala 66:30:@3196.4]
  wire  _T_6001; // @[OneHot.scala 66:30:@3197.4]
  wire  _T_6002; // @[OneHot.scala 66:30:@3198.4]
  wire  _T_6003; // @[OneHot.scala 66:30:@3199.4]
  wire  _T_6004; // @[OneHot.scala 66:30:@3200.4]
  wire  _T_6005; // @[OneHot.scala 66:30:@3201.4]
  wire  _T_6006; // @[OneHot.scala 66:30:@3202.4]
  wire  _T_6007; // @[OneHot.scala 66:30:@3203.4]
  wire  _T_6008; // @[OneHot.scala 66:30:@3204.4]
  wire  _T_6009; // @[OneHot.scala 66:30:@3205.4]
  wire  _T_6010; // @[OneHot.scala 66:30:@3206.4]
  wire [15:0] _T_6051; // @[Mux.scala 31:69:@3224.4]
  wire [15:0] _T_6052; // @[Mux.scala 31:69:@3225.4]
  wire [15:0] _T_6053; // @[Mux.scala 31:69:@3226.4]
  wire [15:0] _T_6054; // @[Mux.scala 31:69:@3227.4]
  wire [15:0] _T_6055; // @[Mux.scala 31:69:@3228.4]
  wire [15:0] _T_6056; // @[Mux.scala 31:69:@3229.4]
  wire [15:0] _T_6057; // @[Mux.scala 31:69:@3230.4]
  wire [15:0] _T_6058; // @[Mux.scala 31:69:@3231.4]
  wire [15:0] _T_6059; // @[Mux.scala 31:69:@3232.4]
  wire [15:0] _T_6060; // @[Mux.scala 31:69:@3233.4]
  wire [15:0] _T_6061; // @[Mux.scala 31:69:@3234.4]
  wire [15:0] _T_6062; // @[Mux.scala 31:69:@3235.4]
  wire [15:0] _T_6063; // @[Mux.scala 31:69:@3236.4]
  wire [15:0] _T_6064; // @[Mux.scala 31:69:@3237.4]
  wire [15:0] _T_6065; // @[Mux.scala 31:69:@3238.4]
  wire [15:0] _T_6066; // @[Mux.scala 31:69:@3239.4]
  wire  _T_6067; // @[OneHot.scala 66:30:@3240.4]
  wire  _T_6068; // @[OneHot.scala 66:30:@3241.4]
  wire  _T_6069; // @[OneHot.scala 66:30:@3242.4]
  wire  _T_6070; // @[OneHot.scala 66:30:@3243.4]
  wire  _T_6071; // @[OneHot.scala 66:30:@3244.4]
  wire  _T_6072; // @[OneHot.scala 66:30:@3245.4]
  wire  _T_6073; // @[OneHot.scala 66:30:@3246.4]
  wire  _T_6074; // @[OneHot.scala 66:30:@3247.4]
  wire  _T_6075; // @[OneHot.scala 66:30:@3248.4]
  wire  _T_6076; // @[OneHot.scala 66:30:@3249.4]
  wire  _T_6077; // @[OneHot.scala 66:30:@3250.4]
  wire  _T_6078; // @[OneHot.scala 66:30:@3251.4]
  wire  _T_6079; // @[OneHot.scala 66:30:@3252.4]
  wire  _T_6080; // @[OneHot.scala 66:30:@3253.4]
  wire  _T_6081; // @[OneHot.scala 66:30:@3254.4]
  wire  _T_6082; // @[OneHot.scala 66:30:@3255.4]
  wire [15:0] _T_6123; // @[Mux.scala 31:69:@3273.4]
  wire [15:0] _T_6124; // @[Mux.scala 31:69:@3274.4]
  wire [15:0] _T_6125; // @[Mux.scala 31:69:@3275.4]
  wire [15:0] _T_6126; // @[Mux.scala 31:69:@3276.4]
  wire [15:0] _T_6127; // @[Mux.scala 31:69:@3277.4]
  wire [15:0] _T_6128; // @[Mux.scala 31:69:@3278.4]
  wire [15:0] _T_6129; // @[Mux.scala 31:69:@3279.4]
  wire [15:0] _T_6130; // @[Mux.scala 31:69:@3280.4]
  wire [15:0] _T_6131; // @[Mux.scala 31:69:@3281.4]
  wire [15:0] _T_6132; // @[Mux.scala 31:69:@3282.4]
  wire [15:0] _T_6133; // @[Mux.scala 31:69:@3283.4]
  wire [15:0] _T_6134; // @[Mux.scala 31:69:@3284.4]
  wire [15:0] _T_6135; // @[Mux.scala 31:69:@3285.4]
  wire [15:0] _T_6136; // @[Mux.scala 31:69:@3286.4]
  wire [15:0] _T_6137; // @[Mux.scala 31:69:@3287.4]
  wire [15:0] _T_6138; // @[Mux.scala 31:69:@3288.4]
  wire  _T_6139; // @[OneHot.scala 66:30:@3289.4]
  wire  _T_6140; // @[OneHot.scala 66:30:@3290.4]
  wire  _T_6141; // @[OneHot.scala 66:30:@3291.4]
  wire  _T_6142; // @[OneHot.scala 66:30:@3292.4]
  wire  _T_6143; // @[OneHot.scala 66:30:@3293.4]
  wire  _T_6144; // @[OneHot.scala 66:30:@3294.4]
  wire  _T_6145; // @[OneHot.scala 66:30:@3295.4]
  wire  _T_6146; // @[OneHot.scala 66:30:@3296.4]
  wire  _T_6147; // @[OneHot.scala 66:30:@3297.4]
  wire  _T_6148; // @[OneHot.scala 66:30:@3298.4]
  wire  _T_6149; // @[OneHot.scala 66:30:@3299.4]
  wire  _T_6150; // @[OneHot.scala 66:30:@3300.4]
  wire  _T_6151; // @[OneHot.scala 66:30:@3301.4]
  wire  _T_6152; // @[OneHot.scala 66:30:@3302.4]
  wire  _T_6153; // @[OneHot.scala 66:30:@3303.4]
  wire  _T_6154; // @[OneHot.scala 66:30:@3304.4]
  wire [15:0] _T_6195; // @[Mux.scala 31:69:@3322.4]
  wire [15:0] _T_6196; // @[Mux.scala 31:69:@3323.4]
  wire [15:0] _T_6197; // @[Mux.scala 31:69:@3324.4]
  wire [15:0] _T_6198; // @[Mux.scala 31:69:@3325.4]
  wire [15:0] _T_6199; // @[Mux.scala 31:69:@3326.4]
  wire [15:0] _T_6200; // @[Mux.scala 31:69:@3327.4]
  wire [15:0] _T_6201; // @[Mux.scala 31:69:@3328.4]
  wire [15:0] _T_6202; // @[Mux.scala 31:69:@3329.4]
  wire [15:0] _T_6203; // @[Mux.scala 31:69:@3330.4]
  wire [15:0] _T_6204; // @[Mux.scala 31:69:@3331.4]
  wire [15:0] _T_6205; // @[Mux.scala 31:69:@3332.4]
  wire [15:0] _T_6206; // @[Mux.scala 31:69:@3333.4]
  wire [15:0] _T_6207; // @[Mux.scala 31:69:@3334.4]
  wire [15:0] _T_6208; // @[Mux.scala 31:69:@3335.4]
  wire [15:0] _T_6209; // @[Mux.scala 31:69:@3336.4]
  wire [15:0] _T_6210; // @[Mux.scala 31:69:@3337.4]
  wire  _T_6211; // @[OneHot.scala 66:30:@3338.4]
  wire  _T_6212; // @[OneHot.scala 66:30:@3339.4]
  wire  _T_6213; // @[OneHot.scala 66:30:@3340.4]
  wire  _T_6214; // @[OneHot.scala 66:30:@3341.4]
  wire  _T_6215; // @[OneHot.scala 66:30:@3342.4]
  wire  _T_6216; // @[OneHot.scala 66:30:@3343.4]
  wire  _T_6217; // @[OneHot.scala 66:30:@3344.4]
  wire  _T_6218; // @[OneHot.scala 66:30:@3345.4]
  wire  _T_6219; // @[OneHot.scala 66:30:@3346.4]
  wire  _T_6220; // @[OneHot.scala 66:30:@3347.4]
  wire  _T_6221; // @[OneHot.scala 66:30:@3348.4]
  wire  _T_6222; // @[OneHot.scala 66:30:@3349.4]
  wire  _T_6223; // @[OneHot.scala 66:30:@3350.4]
  wire  _T_6224; // @[OneHot.scala 66:30:@3351.4]
  wire  _T_6225; // @[OneHot.scala 66:30:@3352.4]
  wire  _T_6226; // @[OneHot.scala 66:30:@3353.4]
  wire [15:0] _T_6267; // @[Mux.scala 31:69:@3371.4]
  wire [15:0] _T_6268; // @[Mux.scala 31:69:@3372.4]
  wire [15:0] _T_6269; // @[Mux.scala 31:69:@3373.4]
  wire [15:0] _T_6270; // @[Mux.scala 31:69:@3374.4]
  wire [15:0] _T_6271; // @[Mux.scala 31:69:@3375.4]
  wire [15:0] _T_6272; // @[Mux.scala 31:69:@3376.4]
  wire [15:0] _T_6273; // @[Mux.scala 31:69:@3377.4]
  wire [15:0] _T_6274; // @[Mux.scala 31:69:@3378.4]
  wire [15:0] _T_6275; // @[Mux.scala 31:69:@3379.4]
  wire [15:0] _T_6276; // @[Mux.scala 31:69:@3380.4]
  wire [15:0] _T_6277; // @[Mux.scala 31:69:@3381.4]
  wire [15:0] _T_6278; // @[Mux.scala 31:69:@3382.4]
  wire [15:0] _T_6279; // @[Mux.scala 31:69:@3383.4]
  wire [15:0] _T_6280; // @[Mux.scala 31:69:@3384.4]
  wire [15:0] _T_6281; // @[Mux.scala 31:69:@3385.4]
  wire [15:0] _T_6282; // @[Mux.scala 31:69:@3386.4]
  wire  _T_6283; // @[OneHot.scala 66:30:@3387.4]
  wire  _T_6284; // @[OneHot.scala 66:30:@3388.4]
  wire  _T_6285; // @[OneHot.scala 66:30:@3389.4]
  wire  _T_6286; // @[OneHot.scala 66:30:@3390.4]
  wire  _T_6287; // @[OneHot.scala 66:30:@3391.4]
  wire  _T_6288; // @[OneHot.scala 66:30:@3392.4]
  wire  _T_6289; // @[OneHot.scala 66:30:@3393.4]
  wire  _T_6290; // @[OneHot.scala 66:30:@3394.4]
  wire  _T_6291; // @[OneHot.scala 66:30:@3395.4]
  wire  _T_6292; // @[OneHot.scala 66:30:@3396.4]
  wire  _T_6293; // @[OneHot.scala 66:30:@3397.4]
  wire  _T_6294; // @[OneHot.scala 66:30:@3398.4]
  wire  _T_6295; // @[OneHot.scala 66:30:@3399.4]
  wire  _T_6296; // @[OneHot.scala 66:30:@3400.4]
  wire  _T_6297; // @[OneHot.scala 66:30:@3401.4]
  wire  _T_6298; // @[OneHot.scala 66:30:@3402.4]
  wire [15:0] _T_6339; // @[Mux.scala 31:69:@3420.4]
  wire [15:0] _T_6340; // @[Mux.scala 31:69:@3421.4]
  wire [15:0] _T_6341; // @[Mux.scala 31:69:@3422.4]
  wire [15:0] _T_6342; // @[Mux.scala 31:69:@3423.4]
  wire [15:0] _T_6343; // @[Mux.scala 31:69:@3424.4]
  wire [15:0] _T_6344; // @[Mux.scala 31:69:@3425.4]
  wire [15:0] _T_6345; // @[Mux.scala 31:69:@3426.4]
  wire [15:0] _T_6346; // @[Mux.scala 31:69:@3427.4]
  wire [15:0] _T_6347; // @[Mux.scala 31:69:@3428.4]
  wire [15:0] _T_6348; // @[Mux.scala 31:69:@3429.4]
  wire [15:0] _T_6349; // @[Mux.scala 31:69:@3430.4]
  wire [15:0] _T_6350; // @[Mux.scala 31:69:@3431.4]
  wire [15:0] _T_6351; // @[Mux.scala 31:69:@3432.4]
  wire [15:0] _T_6352; // @[Mux.scala 31:69:@3433.4]
  wire [15:0] _T_6353; // @[Mux.scala 31:69:@3434.4]
  wire [15:0] _T_6354; // @[Mux.scala 31:69:@3435.4]
  wire  _T_6355; // @[OneHot.scala 66:30:@3436.4]
  wire  _T_6356; // @[OneHot.scala 66:30:@3437.4]
  wire  _T_6357; // @[OneHot.scala 66:30:@3438.4]
  wire  _T_6358; // @[OneHot.scala 66:30:@3439.4]
  wire  _T_6359; // @[OneHot.scala 66:30:@3440.4]
  wire  _T_6360; // @[OneHot.scala 66:30:@3441.4]
  wire  _T_6361; // @[OneHot.scala 66:30:@3442.4]
  wire  _T_6362; // @[OneHot.scala 66:30:@3443.4]
  wire  _T_6363; // @[OneHot.scala 66:30:@3444.4]
  wire  _T_6364; // @[OneHot.scala 66:30:@3445.4]
  wire  _T_6365; // @[OneHot.scala 66:30:@3446.4]
  wire  _T_6366; // @[OneHot.scala 66:30:@3447.4]
  wire  _T_6367; // @[OneHot.scala 66:30:@3448.4]
  wire  _T_6368; // @[OneHot.scala 66:30:@3449.4]
  wire  _T_6369; // @[OneHot.scala 66:30:@3450.4]
  wire  _T_6370; // @[OneHot.scala 66:30:@3451.4]
  wire [15:0] _T_6411; // @[Mux.scala 31:69:@3469.4]
  wire [15:0] _T_6412; // @[Mux.scala 31:69:@3470.4]
  wire [15:0] _T_6413; // @[Mux.scala 31:69:@3471.4]
  wire [15:0] _T_6414; // @[Mux.scala 31:69:@3472.4]
  wire [15:0] _T_6415; // @[Mux.scala 31:69:@3473.4]
  wire [15:0] _T_6416; // @[Mux.scala 31:69:@3474.4]
  wire [15:0] _T_6417; // @[Mux.scala 31:69:@3475.4]
  wire [15:0] _T_6418; // @[Mux.scala 31:69:@3476.4]
  wire [15:0] _T_6419; // @[Mux.scala 31:69:@3477.4]
  wire [15:0] _T_6420; // @[Mux.scala 31:69:@3478.4]
  wire [15:0] _T_6421; // @[Mux.scala 31:69:@3479.4]
  wire [15:0] _T_6422; // @[Mux.scala 31:69:@3480.4]
  wire [15:0] _T_6423; // @[Mux.scala 31:69:@3481.4]
  wire [15:0] _T_6424; // @[Mux.scala 31:69:@3482.4]
  wire [15:0] _T_6425; // @[Mux.scala 31:69:@3483.4]
  wire [15:0] _T_6426; // @[Mux.scala 31:69:@3484.4]
  wire  _T_6427; // @[OneHot.scala 66:30:@3485.4]
  wire  _T_6428; // @[OneHot.scala 66:30:@3486.4]
  wire  _T_6429; // @[OneHot.scala 66:30:@3487.4]
  wire  _T_6430; // @[OneHot.scala 66:30:@3488.4]
  wire  _T_6431; // @[OneHot.scala 66:30:@3489.4]
  wire  _T_6432; // @[OneHot.scala 66:30:@3490.4]
  wire  _T_6433; // @[OneHot.scala 66:30:@3491.4]
  wire  _T_6434; // @[OneHot.scala 66:30:@3492.4]
  wire  _T_6435; // @[OneHot.scala 66:30:@3493.4]
  wire  _T_6436; // @[OneHot.scala 66:30:@3494.4]
  wire  _T_6437; // @[OneHot.scala 66:30:@3495.4]
  wire  _T_6438; // @[OneHot.scala 66:30:@3496.4]
  wire  _T_6439; // @[OneHot.scala 66:30:@3497.4]
  wire  _T_6440; // @[OneHot.scala 66:30:@3498.4]
  wire  _T_6441; // @[OneHot.scala 66:30:@3499.4]
  wire  _T_6442; // @[OneHot.scala 66:30:@3500.4]
  wire [15:0] _T_6483; // @[Mux.scala 31:69:@3518.4]
  wire [15:0] _T_6484; // @[Mux.scala 31:69:@3519.4]
  wire [15:0] _T_6485; // @[Mux.scala 31:69:@3520.4]
  wire [15:0] _T_6486; // @[Mux.scala 31:69:@3521.4]
  wire [15:0] _T_6487; // @[Mux.scala 31:69:@3522.4]
  wire [15:0] _T_6488; // @[Mux.scala 31:69:@3523.4]
  wire [15:0] _T_6489; // @[Mux.scala 31:69:@3524.4]
  wire [15:0] _T_6490; // @[Mux.scala 31:69:@3525.4]
  wire [15:0] _T_6491; // @[Mux.scala 31:69:@3526.4]
  wire [15:0] _T_6492; // @[Mux.scala 31:69:@3527.4]
  wire [15:0] _T_6493; // @[Mux.scala 31:69:@3528.4]
  wire [15:0] _T_6494; // @[Mux.scala 31:69:@3529.4]
  wire [15:0] _T_6495; // @[Mux.scala 31:69:@3530.4]
  wire [15:0] _T_6496; // @[Mux.scala 31:69:@3531.4]
  wire [15:0] _T_6497; // @[Mux.scala 31:69:@3532.4]
  wire [15:0] _T_6498; // @[Mux.scala 31:69:@3533.4]
  wire  _T_6499; // @[OneHot.scala 66:30:@3534.4]
  wire  _T_6500; // @[OneHot.scala 66:30:@3535.4]
  wire  _T_6501; // @[OneHot.scala 66:30:@3536.4]
  wire  _T_6502; // @[OneHot.scala 66:30:@3537.4]
  wire  _T_6503; // @[OneHot.scala 66:30:@3538.4]
  wire  _T_6504; // @[OneHot.scala 66:30:@3539.4]
  wire  _T_6505; // @[OneHot.scala 66:30:@3540.4]
  wire  _T_6506; // @[OneHot.scala 66:30:@3541.4]
  wire  _T_6507; // @[OneHot.scala 66:30:@3542.4]
  wire  _T_6508; // @[OneHot.scala 66:30:@3543.4]
  wire  _T_6509; // @[OneHot.scala 66:30:@3544.4]
  wire  _T_6510; // @[OneHot.scala 66:30:@3545.4]
  wire  _T_6511; // @[OneHot.scala 66:30:@3546.4]
  wire  _T_6512; // @[OneHot.scala 66:30:@3547.4]
  wire  _T_6513; // @[OneHot.scala 66:30:@3548.4]
  wire  _T_6514; // @[OneHot.scala 66:30:@3549.4]
  wire [15:0] _T_6555; // @[Mux.scala 31:69:@3567.4]
  wire [15:0] _T_6556; // @[Mux.scala 31:69:@3568.4]
  wire [15:0] _T_6557; // @[Mux.scala 31:69:@3569.4]
  wire [15:0] _T_6558; // @[Mux.scala 31:69:@3570.4]
  wire [15:0] _T_6559; // @[Mux.scala 31:69:@3571.4]
  wire [15:0] _T_6560; // @[Mux.scala 31:69:@3572.4]
  wire [15:0] _T_6561; // @[Mux.scala 31:69:@3573.4]
  wire [15:0] _T_6562; // @[Mux.scala 31:69:@3574.4]
  wire [15:0] _T_6563; // @[Mux.scala 31:69:@3575.4]
  wire [15:0] _T_6564; // @[Mux.scala 31:69:@3576.4]
  wire [15:0] _T_6565; // @[Mux.scala 31:69:@3577.4]
  wire [15:0] _T_6566; // @[Mux.scala 31:69:@3578.4]
  wire [15:0] _T_6567; // @[Mux.scala 31:69:@3579.4]
  wire [15:0] _T_6568; // @[Mux.scala 31:69:@3580.4]
  wire [15:0] _T_6569; // @[Mux.scala 31:69:@3581.4]
  wire [15:0] _T_6570; // @[Mux.scala 31:69:@3582.4]
  wire  _T_6571; // @[OneHot.scala 66:30:@3583.4]
  wire  _T_6572; // @[OneHot.scala 66:30:@3584.4]
  wire  _T_6573; // @[OneHot.scala 66:30:@3585.4]
  wire  _T_6574; // @[OneHot.scala 66:30:@3586.4]
  wire  _T_6575; // @[OneHot.scala 66:30:@3587.4]
  wire  _T_6576; // @[OneHot.scala 66:30:@3588.4]
  wire  _T_6577; // @[OneHot.scala 66:30:@3589.4]
  wire  _T_6578; // @[OneHot.scala 66:30:@3590.4]
  wire  _T_6579; // @[OneHot.scala 66:30:@3591.4]
  wire  _T_6580; // @[OneHot.scala 66:30:@3592.4]
  wire  _T_6581; // @[OneHot.scala 66:30:@3593.4]
  wire  _T_6582; // @[OneHot.scala 66:30:@3594.4]
  wire  _T_6583; // @[OneHot.scala 66:30:@3595.4]
  wire  _T_6584; // @[OneHot.scala 66:30:@3596.4]
  wire  _T_6585; // @[OneHot.scala 66:30:@3597.4]
  wire  _T_6586; // @[OneHot.scala 66:30:@3598.4]
  wire [15:0] _T_6627; // @[Mux.scala 31:69:@3616.4]
  wire [15:0] _T_6628; // @[Mux.scala 31:69:@3617.4]
  wire [15:0] _T_6629; // @[Mux.scala 31:69:@3618.4]
  wire [15:0] _T_6630; // @[Mux.scala 31:69:@3619.4]
  wire [15:0] _T_6631; // @[Mux.scala 31:69:@3620.4]
  wire [15:0] _T_6632; // @[Mux.scala 31:69:@3621.4]
  wire [15:0] _T_6633; // @[Mux.scala 31:69:@3622.4]
  wire [15:0] _T_6634; // @[Mux.scala 31:69:@3623.4]
  wire [15:0] _T_6635; // @[Mux.scala 31:69:@3624.4]
  wire [15:0] _T_6636; // @[Mux.scala 31:69:@3625.4]
  wire [15:0] _T_6637; // @[Mux.scala 31:69:@3626.4]
  wire [15:0] _T_6638; // @[Mux.scala 31:69:@3627.4]
  wire [15:0] _T_6639; // @[Mux.scala 31:69:@3628.4]
  wire [15:0] _T_6640; // @[Mux.scala 31:69:@3629.4]
  wire [15:0] _T_6641; // @[Mux.scala 31:69:@3630.4]
  wire [15:0] _T_6642; // @[Mux.scala 31:69:@3631.4]
  wire  _T_6643; // @[OneHot.scala 66:30:@3632.4]
  wire  _T_6644; // @[OneHot.scala 66:30:@3633.4]
  wire  _T_6645; // @[OneHot.scala 66:30:@3634.4]
  wire  _T_6646; // @[OneHot.scala 66:30:@3635.4]
  wire  _T_6647; // @[OneHot.scala 66:30:@3636.4]
  wire  _T_6648; // @[OneHot.scala 66:30:@3637.4]
  wire  _T_6649; // @[OneHot.scala 66:30:@3638.4]
  wire  _T_6650; // @[OneHot.scala 66:30:@3639.4]
  wire  _T_6651; // @[OneHot.scala 66:30:@3640.4]
  wire  _T_6652; // @[OneHot.scala 66:30:@3641.4]
  wire  _T_6653; // @[OneHot.scala 66:30:@3642.4]
  wire  _T_6654; // @[OneHot.scala 66:30:@3643.4]
  wire  _T_6655; // @[OneHot.scala 66:30:@3644.4]
  wire  _T_6656; // @[OneHot.scala 66:30:@3645.4]
  wire  _T_6657; // @[OneHot.scala 66:30:@3646.4]
  wire  _T_6658; // @[OneHot.scala 66:30:@3647.4]
  wire [15:0] _T_6699; // @[Mux.scala 31:69:@3665.4]
  wire [15:0] _T_6700; // @[Mux.scala 31:69:@3666.4]
  wire [15:0] _T_6701; // @[Mux.scala 31:69:@3667.4]
  wire [15:0] _T_6702; // @[Mux.scala 31:69:@3668.4]
  wire [15:0] _T_6703; // @[Mux.scala 31:69:@3669.4]
  wire [15:0] _T_6704; // @[Mux.scala 31:69:@3670.4]
  wire [15:0] _T_6705; // @[Mux.scala 31:69:@3671.4]
  wire [15:0] _T_6706; // @[Mux.scala 31:69:@3672.4]
  wire [15:0] _T_6707; // @[Mux.scala 31:69:@3673.4]
  wire [15:0] _T_6708; // @[Mux.scala 31:69:@3674.4]
  wire [15:0] _T_6709; // @[Mux.scala 31:69:@3675.4]
  wire [15:0] _T_6710; // @[Mux.scala 31:69:@3676.4]
  wire [15:0] _T_6711; // @[Mux.scala 31:69:@3677.4]
  wire [15:0] _T_6712; // @[Mux.scala 31:69:@3678.4]
  wire [15:0] _T_6713; // @[Mux.scala 31:69:@3679.4]
  wire [15:0] _T_6714; // @[Mux.scala 31:69:@3680.4]
  wire  _T_6715; // @[OneHot.scala 66:30:@3681.4]
  wire  _T_6716; // @[OneHot.scala 66:30:@3682.4]
  wire  _T_6717; // @[OneHot.scala 66:30:@3683.4]
  wire  _T_6718; // @[OneHot.scala 66:30:@3684.4]
  wire  _T_6719; // @[OneHot.scala 66:30:@3685.4]
  wire  _T_6720; // @[OneHot.scala 66:30:@3686.4]
  wire  _T_6721; // @[OneHot.scala 66:30:@3687.4]
  wire  _T_6722; // @[OneHot.scala 66:30:@3688.4]
  wire  _T_6723; // @[OneHot.scala 66:30:@3689.4]
  wire  _T_6724; // @[OneHot.scala 66:30:@3690.4]
  wire  _T_6725; // @[OneHot.scala 66:30:@3691.4]
  wire  _T_6726; // @[OneHot.scala 66:30:@3692.4]
  wire  _T_6727; // @[OneHot.scala 66:30:@3693.4]
  wire  _T_6728; // @[OneHot.scala 66:30:@3694.4]
  wire  _T_6729; // @[OneHot.scala 66:30:@3695.4]
  wire  _T_6730; // @[OneHot.scala 66:30:@3696.4]
  wire [15:0] _T_6771; // @[Mux.scala 31:69:@3714.4]
  wire [15:0] _T_6772; // @[Mux.scala 31:69:@3715.4]
  wire [15:0] _T_6773; // @[Mux.scala 31:69:@3716.4]
  wire [15:0] _T_6774; // @[Mux.scala 31:69:@3717.4]
  wire [15:0] _T_6775; // @[Mux.scala 31:69:@3718.4]
  wire [15:0] _T_6776; // @[Mux.scala 31:69:@3719.4]
  wire [15:0] _T_6777; // @[Mux.scala 31:69:@3720.4]
  wire [15:0] _T_6778; // @[Mux.scala 31:69:@3721.4]
  wire [15:0] _T_6779; // @[Mux.scala 31:69:@3722.4]
  wire [15:0] _T_6780; // @[Mux.scala 31:69:@3723.4]
  wire [15:0] _T_6781; // @[Mux.scala 31:69:@3724.4]
  wire [15:0] _T_6782; // @[Mux.scala 31:69:@3725.4]
  wire [15:0] _T_6783; // @[Mux.scala 31:69:@3726.4]
  wire [15:0] _T_6784; // @[Mux.scala 31:69:@3727.4]
  wire [15:0] _T_6785; // @[Mux.scala 31:69:@3728.4]
  wire [15:0] _T_6786; // @[Mux.scala 31:69:@3729.4]
  wire  _T_6787; // @[OneHot.scala 66:30:@3730.4]
  wire  _T_6788; // @[OneHot.scala 66:30:@3731.4]
  wire  _T_6789; // @[OneHot.scala 66:30:@3732.4]
  wire  _T_6790; // @[OneHot.scala 66:30:@3733.4]
  wire  _T_6791; // @[OneHot.scala 66:30:@3734.4]
  wire  _T_6792; // @[OneHot.scala 66:30:@3735.4]
  wire  _T_6793; // @[OneHot.scala 66:30:@3736.4]
  wire  _T_6794; // @[OneHot.scala 66:30:@3737.4]
  wire  _T_6795; // @[OneHot.scala 66:30:@3738.4]
  wire  _T_6796; // @[OneHot.scala 66:30:@3739.4]
  wire  _T_6797; // @[OneHot.scala 66:30:@3740.4]
  wire  _T_6798; // @[OneHot.scala 66:30:@3741.4]
  wire  _T_6799; // @[OneHot.scala 66:30:@3742.4]
  wire  _T_6800; // @[OneHot.scala 66:30:@3743.4]
  wire  _T_6801; // @[OneHot.scala 66:30:@3744.4]
  wire  _T_6802; // @[OneHot.scala 66:30:@3745.4]
  wire [15:0] _T_6843; // @[Mux.scala 31:69:@3763.4]
  wire [15:0] _T_6844; // @[Mux.scala 31:69:@3764.4]
  wire [15:0] _T_6845; // @[Mux.scala 31:69:@3765.4]
  wire [15:0] _T_6846; // @[Mux.scala 31:69:@3766.4]
  wire [15:0] _T_6847; // @[Mux.scala 31:69:@3767.4]
  wire [15:0] _T_6848; // @[Mux.scala 31:69:@3768.4]
  wire [15:0] _T_6849; // @[Mux.scala 31:69:@3769.4]
  wire [15:0] _T_6850; // @[Mux.scala 31:69:@3770.4]
  wire [15:0] _T_6851; // @[Mux.scala 31:69:@3771.4]
  wire [15:0] _T_6852; // @[Mux.scala 31:69:@3772.4]
  wire [15:0] _T_6853; // @[Mux.scala 31:69:@3773.4]
  wire [15:0] _T_6854; // @[Mux.scala 31:69:@3774.4]
  wire [15:0] _T_6855; // @[Mux.scala 31:69:@3775.4]
  wire [15:0] _T_6856; // @[Mux.scala 31:69:@3776.4]
  wire [15:0] _T_6857; // @[Mux.scala 31:69:@3777.4]
  wire [15:0] _T_6858; // @[Mux.scala 31:69:@3778.4]
  wire  _T_6859; // @[OneHot.scala 66:30:@3779.4]
  wire  _T_6860; // @[OneHot.scala 66:30:@3780.4]
  wire  _T_6861; // @[OneHot.scala 66:30:@3781.4]
  wire  _T_6862; // @[OneHot.scala 66:30:@3782.4]
  wire  _T_6863; // @[OneHot.scala 66:30:@3783.4]
  wire  _T_6864; // @[OneHot.scala 66:30:@3784.4]
  wire  _T_6865; // @[OneHot.scala 66:30:@3785.4]
  wire  _T_6866; // @[OneHot.scala 66:30:@3786.4]
  wire  _T_6867; // @[OneHot.scala 66:30:@3787.4]
  wire  _T_6868; // @[OneHot.scala 66:30:@3788.4]
  wire  _T_6869; // @[OneHot.scala 66:30:@3789.4]
  wire  _T_6870; // @[OneHot.scala 66:30:@3790.4]
  wire  _T_6871; // @[OneHot.scala 66:30:@3791.4]
  wire  _T_6872; // @[OneHot.scala 66:30:@3792.4]
  wire  _T_6873; // @[OneHot.scala 66:30:@3793.4]
  wire  _T_6874; // @[OneHot.scala 66:30:@3794.4]
  wire [15:0] _T_6915; // @[Mux.scala 31:69:@3812.4]
  wire [15:0] _T_6916; // @[Mux.scala 31:69:@3813.4]
  wire [15:0] _T_6917; // @[Mux.scala 31:69:@3814.4]
  wire [15:0] _T_6918; // @[Mux.scala 31:69:@3815.4]
  wire [15:0] _T_6919; // @[Mux.scala 31:69:@3816.4]
  wire [15:0] _T_6920; // @[Mux.scala 31:69:@3817.4]
  wire [15:0] _T_6921; // @[Mux.scala 31:69:@3818.4]
  wire [15:0] _T_6922; // @[Mux.scala 31:69:@3819.4]
  wire [15:0] _T_6923; // @[Mux.scala 31:69:@3820.4]
  wire [15:0] _T_6924; // @[Mux.scala 31:69:@3821.4]
  wire [15:0] _T_6925; // @[Mux.scala 31:69:@3822.4]
  wire [15:0] _T_6926; // @[Mux.scala 31:69:@3823.4]
  wire [15:0] _T_6927; // @[Mux.scala 31:69:@3824.4]
  wire [15:0] _T_6928; // @[Mux.scala 31:69:@3825.4]
  wire [15:0] _T_6929; // @[Mux.scala 31:69:@3826.4]
  wire [15:0] _T_6930; // @[Mux.scala 31:69:@3827.4]
  wire  _T_6931; // @[OneHot.scala 66:30:@3828.4]
  wire  _T_6932; // @[OneHot.scala 66:30:@3829.4]
  wire  _T_6933; // @[OneHot.scala 66:30:@3830.4]
  wire  _T_6934; // @[OneHot.scala 66:30:@3831.4]
  wire  _T_6935; // @[OneHot.scala 66:30:@3832.4]
  wire  _T_6936; // @[OneHot.scala 66:30:@3833.4]
  wire  _T_6937; // @[OneHot.scala 66:30:@3834.4]
  wire  _T_6938; // @[OneHot.scala 66:30:@3835.4]
  wire  _T_6939; // @[OneHot.scala 66:30:@3836.4]
  wire  _T_6940; // @[OneHot.scala 66:30:@3837.4]
  wire  _T_6941; // @[OneHot.scala 66:30:@3838.4]
  wire  _T_6942; // @[OneHot.scala 66:30:@3839.4]
  wire  _T_6943; // @[OneHot.scala 66:30:@3840.4]
  wire  _T_6944; // @[OneHot.scala 66:30:@3841.4]
  wire  _T_6945; // @[OneHot.scala 66:30:@3842.4]
  wire  _T_6946; // @[OneHot.scala 66:30:@3843.4]
  wire [15:0] _T_6987; // @[Mux.scala 31:69:@3861.4]
  wire [15:0] _T_6988; // @[Mux.scala 31:69:@3862.4]
  wire [15:0] _T_6989; // @[Mux.scala 31:69:@3863.4]
  wire [15:0] _T_6990; // @[Mux.scala 31:69:@3864.4]
  wire [15:0] _T_6991; // @[Mux.scala 31:69:@3865.4]
  wire [15:0] _T_6992; // @[Mux.scala 31:69:@3866.4]
  wire [15:0] _T_6993; // @[Mux.scala 31:69:@3867.4]
  wire [15:0] _T_6994; // @[Mux.scala 31:69:@3868.4]
  wire [15:0] _T_6995; // @[Mux.scala 31:69:@3869.4]
  wire [15:0] _T_6996; // @[Mux.scala 31:69:@3870.4]
  wire [15:0] _T_6997; // @[Mux.scala 31:69:@3871.4]
  wire [15:0] _T_6998; // @[Mux.scala 31:69:@3872.4]
  wire [15:0] _T_6999; // @[Mux.scala 31:69:@3873.4]
  wire [15:0] _T_7000; // @[Mux.scala 31:69:@3874.4]
  wire [15:0] _T_7001; // @[Mux.scala 31:69:@3875.4]
  wire [15:0] _T_7002; // @[Mux.scala 31:69:@3876.4]
  wire  _T_7003; // @[OneHot.scala 66:30:@3877.4]
  wire  _T_7004; // @[OneHot.scala 66:30:@3878.4]
  wire  _T_7005; // @[OneHot.scala 66:30:@3879.4]
  wire  _T_7006; // @[OneHot.scala 66:30:@3880.4]
  wire  _T_7007; // @[OneHot.scala 66:30:@3881.4]
  wire  _T_7008; // @[OneHot.scala 66:30:@3882.4]
  wire  _T_7009; // @[OneHot.scala 66:30:@3883.4]
  wire  _T_7010; // @[OneHot.scala 66:30:@3884.4]
  wire  _T_7011; // @[OneHot.scala 66:30:@3885.4]
  wire  _T_7012; // @[OneHot.scala 66:30:@3886.4]
  wire  _T_7013; // @[OneHot.scala 66:30:@3887.4]
  wire  _T_7014; // @[OneHot.scala 66:30:@3888.4]
  wire  _T_7015; // @[OneHot.scala 66:30:@3889.4]
  wire  _T_7016; // @[OneHot.scala 66:30:@3890.4]
  wire  _T_7017; // @[OneHot.scala 66:30:@3891.4]
  wire  _T_7018; // @[OneHot.scala 66:30:@3892.4]
  wire [15:0] _T_7059; // @[Mux.scala 31:69:@3910.4]
  wire [15:0] _T_7060; // @[Mux.scala 31:69:@3911.4]
  wire [15:0] _T_7061; // @[Mux.scala 31:69:@3912.4]
  wire [15:0] _T_7062; // @[Mux.scala 31:69:@3913.4]
  wire [15:0] _T_7063; // @[Mux.scala 31:69:@3914.4]
  wire [15:0] _T_7064; // @[Mux.scala 31:69:@3915.4]
  wire [15:0] _T_7065; // @[Mux.scala 31:69:@3916.4]
  wire [15:0] _T_7066; // @[Mux.scala 31:69:@3917.4]
  wire [15:0] _T_7067; // @[Mux.scala 31:69:@3918.4]
  wire [15:0] _T_7068; // @[Mux.scala 31:69:@3919.4]
  wire [15:0] _T_7069; // @[Mux.scala 31:69:@3920.4]
  wire [15:0] _T_7070; // @[Mux.scala 31:69:@3921.4]
  wire [15:0] _T_7071; // @[Mux.scala 31:69:@3922.4]
  wire [15:0] _T_7072; // @[Mux.scala 31:69:@3923.4]
  wire [15:0] _T_7073; // @[Mux.scala 31:69:@3924.4]
  wire [15:0] _T_7074; // @[Mux.scala 31:69:@3925.4]
  wire  _T_7075; // @[OneHot.scala 66:30:@3926.4]
  wire  _T_7076; // @[OneHot.scala 66:30:@3927.4]
  wire  _T_7077; // @[OneHot.scala 66:30:@3928.4]
  wire  _T_7078; // @[OneHot.scala 66:30:@3929.4]
  wire  _T_7079; // @[OneHot.scala 66:30:@3930.4]
  wire  _T_7080; // @[OneHot.scala 66:30:@3931.4]
  wire  _T_7081; // @[OneHot.scala 66:30:@3932.4]
  wire  _T_7082; // @[OneHot.scala 66:30:@3933.4]
  wire  _T_7083; // @[OneHot.scala 66:30:@3934.4]
  wire  _T_7084; // @[OneHot.scala 66:30:@3935.4]
  wire  _T_7085; // @[OneHot.scala 66:30:@3936.4]
  wire  _T_7086; // @[OneHot.scala 66:30:@3937.4]
  wire  _T_7087; // @[OneHot.scala 66:30:@3938.4]
  wire  _T_7088; // @[OneHot.scala 66:30:@3939.4]
  wire  _T_7089; // @[OneHot.scala 66:30:@3940.4]
  wire  _T_7090; // @[OneHot.scala 66:30:@3941.4]
  wire [7:0] _T_7155; // @[Mux.scala 19:72:@3965.4]
  wire [15:0] _T_7163; // @[Mux.scala 19:72:@3973.4]
  wire [15:0] _T_7165; // @[Mux.scala 19:72:@3974.4]
  wire [7:0] _T_7172; // @[Mux.scala 19:72:@3981.4]
  wire [15:0] _T_7180; // @[Mux.scala 19:72:@3989.4]
  wire [15:0] _T_7182; // @[Mux.scala 19:72:@3990.4]
  wire [7:0] _T_7189; // @[Mux.scala 19:72:@3997.4]
  wire [15:0] _T_7197; // @[Mux.scala 19:72:@4005.4]
  wire [15:0] _T_7199; // @[Mux.scala 19:72:@4006.4]
  wire [7:0] _T_7206; // @[Mux.scala 19:72:@4013.4]
  wire [15:0] _T_7214; // @[Mux.scala 19:72:@4021.4]
  wire [15:0] _T_7216; // @[Mux.scala 19:72:@4022.4]
  wire [7:0] _T_7223; // @[Mux.scala 19:72:@4029.4]
  wire [15:0] _T_7231; // @[Mux.scala 19:72:@4037.4]
  wire [15:0] _T_7233; // @[Mux.scala 19:72:@4038.4]
  wire [7:0] _T_7240; // @[Mux.scala 19:72:@4045.4]
  wire [15:0] _T_7248; // @[Mux.scala 19:72:@4053.4]
  wire [15:0] _T_7250; // @[Mux.scala 19:72:@4054.4]
  wire [7:0] _T_7257; // @[Mux.scala 19:72:@4061.4]
  wire [15:0] _T_7265; // @[Mux.scala 19:72:@4069.4]
  wire [15:0] _T_7267; // @[Mux.scala 19:72:@4070.4]
  wire [7:0] _T_7274; // @[Mux.scala 19:72:@4077.4]
  wire [15:0] _T_7282; // @[Mux.scala 19:72:@4085.4]
  wire [15:0] _T_7284; // @[Mux.scala 19:72:@4086.4]
  wire [7:0] _T_7291; // @[Mux.scala 19:72:@4093.4]
  wire [15:0] _T_7299; // @[Mux.scala 19:72:@4101.4]
  wire [15:0] _T_7301; // @[Mux.scala 19:72:@4102.4]
  wire [7:0] _T_7308; // @[Mux.scala 19:72:@4109.4]
  wire [15:0] _T_7316; // @[Mux.scala 19:72:@4117.4]
  wire [15:0] _T_7318; // @[Mux.scala 19:72:@4118.4]
  wire [7:0] _T_7325; // @[Mux.scala 19:72:@4125.4]
  wire [15:0] _T_7333; // @[Mux.scala 19:72:@4133.4]
  wire [15:0] _T_7335; // @[Mux.scala 19:72:@4134.4]
  wire [7:0] _T_7342; // @[Mux.scala 19:72:@4141.4]
  wire [15:0] _T_7350; // @[Mux.scala 19:72:@4149.4]
  wire [15:0] _T_7352; // @[Mux.scala 19:72:@4150.4]
  wire [7:0] _T_7359; // @[Mux.scala 19:72:@4157.4]
  wire [15:0] _T_7367; // @[Mux.scala 19:72:@4165.4]
  wire [15:0] _T_7369; // @[Mux.scala 19:72:@4166.4]
  wire [7:0] _T_7376; // @[Mux.scala 19:72:@4173.4]
  wire [15:0] _T_7384; // @[Mux.scala 19:72:@4181.4]
  wire [15:0] _T_7386; // @[Mux.scala 19:72:@4182.4]
  wire [7:0] _T_7393; // @[Mux.scala 19:72:@4189.4]
  wire [15:0] _T_7401; // @[Mux.scala 19:72:@4197.4]
  wire [15:0] _T_7403; // @[Mux.scala 19:72:@4198.4]
  wire [7:0] _T_7410; // @[Mux.scala 19:72:@4205.4]
  wire [15:0] _T_7418; // @[Mux.scala 19:72:@4213.4]
  wire [15:0] _T_7420; // @[Mux.scala 19:72:@4214.4]
  wire [15:0] _T_7421; // @[Mux.scala 19:72:@4215.4]
  wire [15:0] _T_7422; // @[Mux.scala 19:72:@4216.4]
  wire [15:0] _T_7423; // @[Mux.scala 19:72:@4217.4]
  wire [15:0] _T_7424; // @[Mux.scala 19:72:@4218.4]
  wire [15:0] _T_7425; // @[Mux.scala 19:72:@4219.4]
  wire [15:0] _T_7426; // @[Mux.scala 19:72:@4220.4]
  wire [15:0] _T_7427; // @[Mux.scala 19:72:@4221.4]
  wire [15:0] _T_7428; // @[Mux.scala 19:72:@4222.4]
  wire [15:0] _T_7429; // @[Mux.scala 19:72:@4223.4]
  wire [15:0] _T_7430; // @[Mux.scala 19:72:@4224.4]
  wire [15:0] _T_7431; // @[Mux.scala 19:72:@4225.4]
  wire [15:0] _T_7432; // @[Mux.scala 19:72:@4226.4]
  wire [15:0] _T_7433; // @[Mux.scala 19:72:@4227.4]
  wire [15:0] _T_7434; // @[Mux.scala 19:72:@4228.4]
  wire [15:0] _T_7435; // @[Mux.scala 19:72:@4229.4]
  wire  inputDataPriorityPorts_0_0; // @[Mux.scala 19:72:@4233.4]
  wire  inputDataPriorityPorts_0_1; // @[Mux.scala 19:72:@4235.4]
  wire  inputDataPriorityPorts_0_2; // @[Mux.scala 19:72:@4237.4]
  wire  inputDataPriorityPorts_0_3; // @[Mux.scala 19:72:@4239.4]
  wire  inputDataPriorityPorts_0_4; // @[Mux.scala 19:72:@4241.4]
  wire  inputDataPriorityPorts_0_5; // @[Mux.scala 19:72:@4243.4]
  wire  inputDataPriorityPorts_0_6; // @[Mux.scala 19:72:@4245.4]
  wire  inputDataPriorityPorts_0_7; // @[Mux.scala 19:72:@4247.4]
  wire  inputDataPriorityPorts_0_8; // @[Mux.scala 19:72:@4249.4]
  wire  inputDataPriorityPorts_0_9; // @[Mux.scala 19:72:@4251.4]
  wire  inputDataPriorityPorts_0_10; // @[Mux.scala 19:72:@4253.4]
  wire  inputDataPriorityPorts_0_11; // @[Mux.scala 19:72:@4255.4]
  wire  inputDataPriorityPorts_0_12; // @[Mux.scala 19:72:@4257.4]
  wire  inputDataPriorityPorts_0_13; // @[Mux.scala 19:72:@4259.4]
  wire  inputDataPriorityPorts_0_14; // @[Mux.scala 19:72:@4261.4]
  wire  inputDataPriorityPorts_0_15; // @[Mux.scala 19:72:@4263.4]
  wire  _T_7581; // @[StoreQueue.scala 209:52:@4287.6]
  wire  _T_7582; // @[StoreQueue.scala 209:81:@4288.6]
  wire [31:0] _GEN_992; // @[StoreQueue.scala 210:40:@4292.6]
  wire  _GEN_993; // @[StoreQueue.scala 210:40:@4292.6]
  wire  _T_7598; // @[StoreQueue.scala 215:52:@4297.6]
  wire  _T_7599; // @[StoreQueue.scala 215:81:@4298.6]
  wire [31:0] _GEN_994; // @[StoreQueue.scala 216:40:@4302.6]
  wire  _GEN_995; // @[StoreQueue.scala 216:40:@4302.6]
  wire  _GEN_996; // @[StoreQueue.scala 204:35:@4281.4]
  wire  _GEN_997; // @[StoreQueue.scala 204:35:@4281.4]
  wire [31:0] _GEN_998; // @[StoreQueue.scala 204:35:@4281.4]
  wire [31:0] _GEN_999; // @[StoreQueue.scala 204:35:@4281.4]
  wire  _T_7617; // @[StoreQueue.scala 209:52:@4313.6]
  wire  _T_7618; // @[StoreQueue.scala 209:81:@4314.6]
  wire [31:0] _GEN_1000; // @[StoreQueue.scala 210:40:@4318.6]
  wire  _GEN_1001; // @[StoreQueue.scala 210:40:@4318.6]
  wire  _T_7634; // @[StoreQueue.scala 215:52:@4323.6]
  wire  _T_7635; // @[StoreQueue.scala 215:81:@4324.6]
  wire [31:0] _GEN_1002; // @[StoreQueue.scala 216:40:@4328.6]
  wire  _GEN_1003; // @[StoreQueue.scala 216:40:@4328.6]
  wire  _GEN_1004; // @[StoreQueue.scala 204:35:@4307.4]
  wire  _GEN_1005; // @[StoreQueue.scala 204:35:@4307.4]
  wire [31:0] _GEN_1006; // @[StoreQueue.scala 204:35:@4307.4]
  wire [31:0] _GEN_1007; // @[StoreQueue.scala 204:35:@4307.4]
  wire  _T_7653; // @[StoreQueue.scala 209:52:@4339.6]
  wire  _T_7654; // @[StoreQueue.scala 209:81:@4340.6]
  wire [31:0] _GEN_1008; // @[StoreQueue.scala 210:40:@4344.6]
  wire  _GEN_1009; // @[StoreQueue.scala 210:40:@4344.6]
  wire  _T_7670; // @[StoreQueue.scala 215:52:@4349.6]
  wire  _T_7671; // @[StoreQueue.scala 215:81:@4350.6]
  wire [31:0] _GEN_1010; // @[StoreQueue.scala 216:40:@4354.6]
  wire  _GEN_1011; // @[StoreQueue.scala 216:40:@4354.6]
  wire  _GEN_1012; // @[StoreQueue.scala 204:35:@4333.4]
  wire  _GEN_1013; // @[StoreQueue.scala 204:35:@4333.4]
  wire [31:0] _GEN_1014; // @[StoreQueue.scala 204:35:@4333.4]
  wire [31:0] _GEN_1015; // @[StoreQueue.scala 204:35:@4333.4]
  wire  _T_7689; // @[StoreQueue.scala 209:52:@4365.6]
  wire  _T_7690; // @[StoreQueue.scala 209:81:@4366.6]
  wire [31:0] _GEN_1016; // @[StoreQueue.scala 210:40:@4370.6]
  wire  _GEN_1017; // @[StoreQueue.scala 210:40:@4370.6]
  wire  _T_7706; // @[StoreQueue.scala 215:52:@4375.6]
  wire  _T_7707; // @[StoreQueue.scala 215:81:@4376.6]
  wire [31:0] _GEN_1018; // @[StoreQueue.scala 216:40:@4380.6]
  wire  _GEN_1019; // @[StoreQueue.scala 216:40:@4380.6]
  wire  _GEN_1020; // @[StoreQueue.scala 204:35:@4359.4]
  wire  _GEN_1021; // @[StoreQueue.scala 204:35:@4359.4]
  wire [31:0] _GEN_1022; // @[StoreQueue.scala 204:35:@4359.4]
  wire [31:0] _GEN_1023; // @[StoreQueue.scala 204:35:@4359.4]
  wire  _T_7725; // @[StoreQueue.scala 209:52:@4391.6]
  wire  _T_7726; // @[StoreQueue.scala 209:81:@4392.6]
  wire [31:0] _GEN_1024; // @[StoreQueue.scala 210:40:@4396.6]
  wire  _GEN_1025; // @[StoreQueue.scala 210:40:@4396.6]
  wire  _T_7742; // @[StoreQueue.scala 215:52:@4401.6]
  wire  _T_7743; // @[StoreQueue.scala 215:81:@4402.6]
  wire [31:0] _GEN_1026; // @[StoreQueue.scala 216:40:@4406.6]
  wire  _GEN_1027; // @[StoreQueue.scala 216:40:@4406.6]
  wire  _GEN_1028; // @[StoreQueue.scala 204:35:@4385.4]
  wire  _GEN_1029; // @[StoreQueue.scala 204:35:@4385.4]
  wire [31:0] _GEN_1030; // @[StoreQueue.scala 204:35:@4385.4]
  wire [31:0] _GEN_1031; // @[StoreQueue.scala 204:35:@4385.4]
  wire  _T_7761; // @[StoreQueue.scala 209:52:@4417.6]
  wire  _T_7762; // @[StoreQueue.scala 209:81:@4418.6]
  wire [31:0] _GEN_1032; // @[StoreQueue.scala 210:40:@4422.6]
  wire  _GEN_1033; // @[StoreQueue.scala 210:40:@4422.6]
  wire  _T_7778; // @[StoreQueue.scala 215:52:@4427.6]
  wire  _T_7779; // @[StoreQueue.scala 215:81:@4428.6]
  wire [31:0] _GEN_1034; // @[StoreQueue.scala 216:40:@4432.6]
  wire  _GEN_1035; // @[StoreQueue.scala 216:40:@4432.6]
  wire  _GEN_1036; // @[StoreQueue.scala 204:35:@4411.4]
  wire  _GEN_1037; // @[StoreQueue.scala 204:35:@4411.4]
  wire [31:0] _GEN_1038; // @[StoreQueue.scala 204:35:@4411.4]
  wire [31:0] _GEN_1039; // @[StoreQueue.scala 204:35:@4411.4]
  wire  _T_7797; // @[StoreQueue.scala 209:52:@4443.6]
  wire  _T_7798; // @[StoreQueue.scala 209:81:@4444.6]
  wire [31:0] _GEN_1040; // @[StoreQueue.scala 210:40:@4448.6]
  wire  _GEN_1041; // @[StoreQueue.scala 210:40:@4448.6]
  wire  _T_7814; // @[StoreQueue.scala 215:52:@4453.6]
  wire  _T_7815; // @[StoreQueue.scala 215:81:@4454.6]
  wire [31:0] _GEN_1042; // @[StoreQueue.scala 216:40:@4458.6]
  wire  _GEN_1043; // @[StoreQueue.scala 216:40:@4458.6]
  wire  _GEN_1044; // @[StoreQueue.scala 204:35:@4437.4]
  wire  _GEN_1045; // @[StoreQueue.scala 204:35:@4437.4]
  wire [31:0] _GEN_1046; // @[StoreQueue.scala 204:35:@4437.4]
  wire [31:0] _GEN_1047; // @[StoreQueue.scala 204:35:@4437.4]
  wire  _T_7833; // @[StoreQueue.scala 209:52:@4469.6]
  wire  _T_7834; // @[StoreQueue.scala 209:81:@4470.6]
  wire [31:0] _GEN_1048; // @[StoreQueue.scala 210:40:@4474.6]
  wire  _GEN_1049; // @[StoreQueue.scala 210:40:@4474.6]
  wire  _T_7850; // @[StoreQueue.scala 215:52:@4479.6]
  wire  _T_7851; // @[StoreQueue.scala 215:81:@4480.6]
  wire [31:0] _GEN_1050; // @[StoreQueue.scala 216:40:@4484.6]
  wire  _GEN_1051; // @[StoreQueue.scala 216:40:@4484.6]
  wire  _GEN_1052; // @[StoreQueue.scala 204:35:@4463.4]
  wire  _GEN_1053; // @[StoreQueue.scala 204:35:@4463.4]
  wire [31:0] _GEN_1054; // @[StoreQueue.scala 204:35:@4463.4]
  wire [31:0] _GEN_1055; // @[StoreQueue.scala 204:35:@4463.4]
  wire  _T_7869; // @[StoreQueue.scala 209:52:@4495.6]
  wire  _T_7870; // @[StoreQueue.scala 209:81:@4496.6]
  wire [31:0] _GEN_1056; // @[StoreQueue.scala 210:40:@4500.6]
  wire  _GEN_1057; // @[StoreQueue.scala 210:40:@4500.6]
  wire  _T_7886; // @[StoreQueue.scala 215:52:@4505.6]
  wire  _T_7887; // @[StoreQueue.scala 215:81:@4506.6]
  wire [31:0] _GEN_1058; // @[StoreQueue.scala 216:40:@4510.6]
  wire  _GEN_1059; // @[StoreQueue.scala 216:40:@4510.6]
  wire  _GEN_1060; // @[StoreQueue.scala 204:35:@4489.4]
  wire  _GEN_1061; // @[StoreQueue.scala 204:35:@4489.4]
  wire [31:0] _GEN_1062; // @[StoreQueue.scala 204:35:@4489.4]
  wire [31:0] _GEN_1063; // @[StoreQueue.scala 204:35:@4489.4]
  wire  _T_7905; // @[StoreQueue.scala 209:52:@4521.6]
  wire  _T_7906; // @[StoreQueue.scala 209:81:@4522.6]
  wire [31:0] _GEN_1064; // @[StoreQueue.scala 210:40:@4526.6]
  wire  _GEN_1065; // @[StoreQueue.scala 210:40:@4526.6]
  wire  _T_7922; // @[StoreQueue.scala 215:52:@4531.6]
  wire  _T_7923; // @[StoreQueue.scala 215:81:@4532.6]
  wire [31:0] _GEN_1066; // @[StoreQueue.scala 216:40:@4536.6]
  wire  _GEN_1067; // @[StoreQueue.scala 216:40:@4536.6]
  wire  _GEN_1068; // @[StoreQueue.scala 204:35:@4515.4]
  wire  _GEN_1069; // @[StoreQueue.scala 204:35:@4515.4]
  wire [31:0] _GEN_1070; // @[StoreQueue.scala 204:35:@4515.4]
  wire [31:0] _GEN_1071; // @[StoreQueue.scala 204:35:@4515.4]
  wire  _T_7941; // @[StoreQueue.scala 209:52:@4547.6]
  wire  _T_7942; // @[StoreQueue.scala 209:81:@4548.6]
  wire [31:0] _GEN_1072; // @[StoreQueue.scala 210:40:@4552.6]
  wire  _GEN_1073; // @[StoreQueue.scala 210:40:@4552.6]
  wire  _T_7958; // @[StoreQueue.scala 215:52:@4557.6]
  wire  _T_7959; // @[StoreQueue.scala 215:81:@4558.6]
  wire [31:0] _GEN_1074; // @[StoreQueue.scala 216:40:@4562.6]
  wire  _GEN_1075; // @[StoreQueue.scala 216:40:@4562.6]
  wire  _GEN_1076; // @[StoreQueue.scala 204:35:@4541.4]
  wire  _GEN_1077; // @[StoreQueue.scala 204:35:@4541.4]
  wire [31:0] _GEN_1078; // @[StoreQueue.scala 204:35:@4541.4]
  wire [31:0] _GEN_1079; // @[StoreQueue.scala 204:35:@4541.4]
  wire  _T_7977; // @[StoreQueue.scala 209:52:@4573.6]
  wire  _T_7978; // @[StoreQueue.scala 209:81:@4574.6]
  wire [31:0] _GEN_1080; // @[StoreQueue.scala 210:40:@4578.6]
  wire  _GEN_1081; // @[StoreQueue.scala 210:40:@4578.6]
  wire  _T_7994; // @[StoreQueue.scala 215:52:@4583.6]
  wire  _T_7995; // @[StoreQueue.scala 215:81:@4584.6]
  wire [31:0] _GEN_1082; // @[StoreQueue.scala 216:40:@4588.6]
  wire  _GEN_1083; // @[StoreQueue.scala 216:40:@4588.6]
  wire  _GEN_1084; // @[StoreQueue.scala 204:35:@4567.4]
  wire  _GEN_1085; // @[StoreQueue.scala 204:35:@4567.4]
  wire [31:0] _GEN_1086; // @[StoreQueue.scala 204:35:@4567.4]
  wire [31:0] _GEN_1087; // @[StoreQueue.scala 204:35:@4567.4]
  wire  _T_8013; // @[StoreQueue.scala 209:52:@4599.6]
  wire  _T_8014; // @[StoreQueue.scala 209:81:@4600.6]
  wire [31:0] _GEN_1088; // @[StoreQueue.scala 210:40:@4604.6]
  wire  _GEN_1089; // @[StoreQueue.scala 210:40:@4604.6]
  wire  _T_8030; // @[StoreQueue.scala 215:52:@4609.6]
  wire  _T_8031; // @[StoreQueue.scala 215:81:@4610.6]
  wire [31:0] _GEN_1090; // @[StoreQueue.scala 216:40:@4614.6]
  wire  _GEN_1091; // @[StoreQueue.scala 216:40:@4614.6]
  wire  _GEN_1092; // @[StoreQueue.scala 204:35:@4593.4]
  wire  _GEN_1093; // @[StoreQueue.scala 204:35:@4593.4]
  wire [31:0] _GEN_1094; // @[StoreQueue.scala 204:35:@4593.4]
  wire [31:0] _GEN_1095; // @[StoreQueue.scala 204:35:@4593.4]
  wire  _T_8049; // @[StoreQueue.scala 209:52:@4625.6]
  wire  _T_8050; // @[StoreQueue.scala 209:81:@4626.6]
  wire [31:0] _GEN_1096; // @[StoreQueue.scala 210:40:@4630.6]
  wire  _GEN_1097; // @[StoreQueue.scala 210:40:@4630.6]
  wire  _T_8066; // @[StoreQueue.scala 215:52:@4635.6]
  wire  _T_8067; // @[StoreQueue.scala 215:81:@4636.6]
  wire [31:0] _GEN_1098; // @[StoreQueue.scala 216:40:@4640.6]
  wire  _GEN_1099; // @[StoreQueue.scala 216:40:@4640.6]
  wire  _GEN_1100; // @[StoreQueue.scala 204:35:@4619.4]
  wire  _GEN_1101; // @[StoreQueue.scala 204:35:@4619.4]
  wire [31:0] _GEN_1102; // @[StoreQueue.scala 204:35:@4619.4]
  wire [31:0] _GEN_1103; // @[StoreQueue.scala 204:35:@4619.4]
  wire  _T_8085; // @[StoreQueue.scala 209:52:@4651.6]
  wire  _T_8086; // @[StoreQueue.scala 209:81:@4652.6]
  wire [31:0] _GEN_1104; // @[StoreQueue.scala 210:40:@4656.6]
  wire  _GEN_1105; // @[StoreQueue.scala 210:40:@4656.6]
  wire  _T_8102; // @[StoreQueue.scala 215:52:@4661.6]
  wire  _T_8103; // @[StoreQueue.scala 215:81:@4662.6]
  wire [31:0] _GEN_1106; // @[StoreQueue.scala 216:40:@4666.6]
  wire  _GEN_1107; // @[StoreQueue.scala 216:40:@4666.6]
  wire  _GEN_1108; // @[StoreQueue.scala 204:35:@4645.4]
  wire  _GEN_1109; // @[StoreQueue.scala 204:35:@4645.4]
  wire [31:0] _GEN_1110; // @[StoreQueue.scala 204:35:@4645.4]
  wire [31:0] _GEN_1111; // @[StoreQueue.scala 204:35:@4645.4]
  wire  _T_8121; // @[StoreQueue.scala 209:52:@4677.6]
  wire  _T_8122; // @[StoreQueue.scala 209:81:@4678.6]
  wire [31:0] _GEN_1112; // @[StoreQueue.scala 210:40:@4682.6]
  wire  _GEN_1113; // @[StoreQueue.scala 210:40:@4682.6]
  wire  _T_8138; // @[StoreQueue.scala 215:52:@4687.6]
  wire  _T_8139; // @[StoreQueue.scala 215:81:@4688.6]
  wire [31:0] _GEN_1114; // @[StoreQueue.scala 216:40:@4692.6]
  wire  _GEN_1115; // @[StoreQueue.scala 216:40:@4692.6]
  wire  _GEN_1116; // @[StoreQueue.scala 204:35:@4671.4]
  wire  _GEN_1117; // @[StoreQueue.scala 204:35:@4671.4]
  wire [31:0] _GEN_1118; // @[StoreQueue.scala 204:35:@4671.4]
  wire [31:0] _GEN_1119; // @[StoreQueue.scala 204:35:@4671.4]
  wire  _T_8153; // @[StoreQueue.scala 229:23:@4697.4]
  wire [4:0] _T_8156; // @[util.scala 10:8:@4699.6]
  wire [4:0] _GEN_64; // @[util.scala 10:14:@4700.6]
  wire [4:0] _T_8157; // @[util.scala 10:14:@4700.6]
  wire [4:0] _GEN_1120; // @[StoreQueue.scala 229:50:@4698.4]
  wire [3:0] _GEN_1234; // @[util.scala 10:8:@4704.6]
  wire [4:0] _T_8159; // @[util.scala 10:8:@4704.6]
  wire [4:0] _GEN_65; // @[util.scala 10:14:@4705.6]
  wire [4:0] _T_8160; // @[util.scala 10:14:@4705.6]
  wire [4:0] _GEN_1121; // @[StoreQueue.scala 233:20:@4703.4]
  wire  _T_8162; // @[StoreQueue.scala 237:84:@4708.4]
  wire  _T_8163; // @[StoreQueue.scala 237:81:@4709.4]
  wire  _T_8165; // @[StoreQueue.scala 237:84:@4710.4]
  wire  _T_8166; // @[StoreQueue.scala 237:81:@4711.4]
  wire  _T_8168; // @[StoreQueue.scala 237:84:@4712.4]
  wire  _T_8169; // @[StoreQueue.scala 237:81:@4713.4]
  wire  _T_8171; // @[StoreQueue.scala 237:84:@4714.4]
  wire  _T_8172; // @[StoreQueue.scala 237:81:@4715.4]
  wire  _T_8174; // @[StoreQueue.scala 237:84:@4716.4]
  wire  _T_8175; // @[StoreQueue.scala 237:81:@4717.4]
  wire  _T_8177; // @[StoreQueue.scala 237:84:@4718.4]
  wire  _T_8178; // @[StoreQueue.scala 237:81:@4719.4]
  wire  _T_8180; // @[StoreQueue.scala 237:84:@4720.4]
  wire  _T_8181; // @[StoreQueue.scala 237:81:@4721.4]
  wire  _T_8183; // @[StoreQueue.scala 237:84:@4722.4]
  wire  _T_8184; // @[StoreQueue.scala 237:81:@4723.4]
  wire  _T_8186; // @[StoreQueue.scala 237:84:@4724.4]
  wire  _T_8187; // @[StoreQueue.scala 237:81:@4725.4]
  wire  _T_8189; // @[StoreQueue.scala 237:84:@4726.4]
  wire  _T_8190; // @[StoreQueue.scala 237:81:@4727.4]
  wire  _T_8192; // @[StoreQueue.scala 237:84:@4728.4]
  wire  _T_8193; // @[StoreQueue.scala 237:81:@4729.4]
  wire  _T_8195; // @[StoreQueue.scala 237:84:@4730.4]
  wire  _T_8196; // @[StoreQueue.scala 237:81:@4731.4]
  wire  _T_8198; // @[StoreQueue.scala 237:84:@4732.4]
  wire  _T_8199; // @[StoreQueue.scala 237:81:@4733.4]
  wire  _T_8201; // @[StoreQueue.scala 237:84:@4734.4]
  wire  _T_8202; // @[StoreQueue.scala 237:81:@4735.4]
  wire  _T_8204; // @[StoreQueue.scala 237:84:@4736.4]
  wire  _T_8205; // @[StoreQueue.scala 237:81:@4737.4]
  wire  _T_8207; // @[StoreQueue.scala 237:84:@4738.4]
  wire  _T_8208; // @[StoreQueue.scala 237:81:@4739.4]
  wire  _T_8233; // @[StoreQueue.scala 237:98:@4758.4]
  wire  _T_8234; // @[StoreQueue.scala 237:98:@4759.4]
  wire  _T_8235; // @[StoreQueue.scala 237:98:@4760.4]
  wire  _T_8236; // @[StoreQueue.scala 237:98:@4761.4]
  wire  _T_8237; // @[StoreQueue.scala 237:98:@4762.4]
  wire  _T_8238; // @[StoreQueue.scala 237:98:@4763.4]
  wire  _T_8239; // @[StoreQueue.scala 237:98:@4764.4]
  wire  _T_8240; // @[StoreQueue.scala 237:98:@4765.4]
  wire  _T_8241; // @[StoreQueue.scala 237:98:@4766.4]
  wire  _T_8242; // @[StoreQueue.scala 237:98:@4767.4]
  wire  _T_8243; // @[StoreQueue.scala 237:98:@4768.4]
  wire  _T_8244; // @[StoreQueue.scala 237:98:@4769.4]
  wire  _T_8245; // @[StoreQueue.scala 237:98:@4770.4]
  wire  _T_8246; // @[StoreQueue.scala 237:98:@4771.4]
  wire [31:0] _GEN_1123; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1124; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1125; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1126; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1127; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1128; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1129; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1130; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1131; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1132; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1133; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1134; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1135; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1136; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1138 = {{2'd0}, tail}; // @[util.scala 14:20:@173.4]
  assign _T_1596 = 6'h10 - _GEN_1138; // @[util.scala 14:20:@173.4]
  assign _T_1597 = $unsigned(_T_1596); // @[util.scala 14:20:@174.4]
  assign _T_1598 = _T_1597[5:0]; // @[util.scala 14:20:@175.4]
  assign _GEN_0 = _T_1598 % 6'h10; // @[util.scala 14:25:@176.4]
  assign _T_1599 = _GEN_0[4:0]; // @[util.scala 14:25:@176.4]
  assign _GEN_1139 = {{3'd0}, io_bbNumStores}; // @[StoreQueue.scala 70:46:@177.4]
  assign _T_1600 = _T_1599 < _GEN_1139; // @[StoreQueue.scala 70:46:@177.4]
  assign initBits_0 = _T_1600 & io_bbStart; // @[StoreQueue.scala 70:64:@178.4]
  assign _T_1605 = 6'h11 - _GEN_1138; // @[util.scala 14:20:@180.4]
  assign _T_1606 = $unsigned(_T_1605); // @[util.scala 14:20:@181.4]
  assign _T_1607 = _T_1606[5:0]; // @[util.scala 14:20:@182.4]
  assign _GEN_16 = _T_1607 % 6'h10; // @[util.scala 14:25:@183.4]
  assign _T_1608 = _GEN_16[4:0]; // @[util.scala 14:25:@183.4]
  assign _T_1609 = _T_1608 < _GEN_1139; // @[StoreQueue.scala 70:46:@184.4]
  assign initBits_1 = _T_1609 & io_bbStart; // @[StoreQueue.scala 70:64:@185.4]
  assign _T_1614 = 6'h12 - _GEN_1138; // @[util.scala 14:20:@187.4]
  assign _T_1615 = $unsigned(_T_1614); // @[util.scala 14:20:@188.4]
  assign _T_1616 = _T_1615[5:0]; // @[util.scala 14:20:@189.4]
  assign _GEN_17 = _T_1616 % 6'h10; // @[util.scala 14:25:@190.4]
  assign _T_1617 = _GEN_17[4:0]; // @[util.scala 14:25:@190.4]
  assign _T_1618 = _T_1617 < _GEN_1139; // @[StoreQueue.scala 70:46:@191.4]
  assign initBits_2 = _T_1618 & io_bbStart; // @[StoreQueue.scala 70:64:@192.4]
  assign _T_1623 = 6'h13 - _GEN_1138; // @[util.scala 14:20:@194.4]
  assign _T_1624 = $unsigned(_T_1623); // @[util.scala 14:20:@195.4]
  assign _T_1625 = _T_1624[5:0]; // @[util.scala 14:20:@196.4]
  assign _GEN_18 = _T_1625 % 6'h10; // @[util.scala 14:25:@197.4]
  assign _T_1626 = _GEN_18[4:0]; // @[util.scala 14:25:@197.4]
  assign _T_1627 = _T_1626 < _GEN_1139; // @[StoreQueue.scala 70:46:@198.4]
  assign initBits_3 = _T_1627 & io_bbStart; // @[StoreQueue.scala 70:64:@199.4]
  assign _T_1632 = 6'h14 - _GEN_1138; // @[util.scala 14:20:@201.4]
  assign _T_1633 = $unsigned(_T_1632); // @[util.scala 14:20:@202.4]
  assign _T_1634 = _T_1633[5:0]; // @[util.scala 14:20:@203.4]
  assign _GEN_19 = _T_1634 % 6'h10; // @[util.scala 14:25:@204.4]
  assign _T_1635 = _GEN_19[4:0]; // @[util.scala 14:25:@204.4]
  assign _T_1636 = _T_1635 < _GEN_1139; // @[StoreQueue.scala 70:46:@205.4]
  assign initBits_4 = _T_1636 & io_bbStart; // @[StoreQueue.scala 70:64:@206.4]
  assign _T_1641 = 6'h15 - _GEN_1138; // @[util.scala 14:20:@208.4]
  assign _T_1642 = $unsigned(_T_1641); // @[util.scala 14:20:@209.4]
  assign _T_1643 = _T_1642[5:0]; // @[util.scala 14:20:@210.4]
  assign _GEN_20 = _T_1643 % 6'h10; // @[util.scala 14:25:@211.4]
  assign _T_1644 = _GEN_20[4:0]; // @[util.scala 14:25:@211.4]
  assign _T_1645 = _T_1644 < _GEN_1139; // @[StoreQueue.scala 70:46:@212.4]
  assign initBits_5 = _T_1645 & io_bbStart; // @[StoreQueue.scala 70:64:@213.4]
  assign _T_1650 = 6'h16 - _GEN_1138; // @[util.scala 14:20:@215.4]
  assign _T_1651 = $unsigned(_T_1650); // @[util.scala 14:20:@216.4]
  assign _T_1652 = _T_1651[5:0]; // @[util.scala 14:20:@217.4]
  assign _GEN_21 = _T_1652 % 6'h10; // @[util.scala 14:25:@218.4]
  assign _T_1653 = _GEN_21[4:0]; // @[util.scala 14:25:@218.4]
  assign _T_1654 = _T_1653 < _GEN_1139; // @[StoreQueue.scala 70:46:@219.4]
  assign initBits_6 = _T_1654 & io_bbStart; // @[StoreQueue.scala 70:64:@220.4]
  assign _T_1659 = 6'h17 - _GEN_1138; // @[util.scala 14:20:@222.4]
  assign _T_1660 = $unsigned(_T_1659); // @[util.scala 14:20:@223.4]
  assign _T_1661 = _T_1660[5:0]; // @[util.scala 14:20:@224.4]
  assign _GEN_22 = _T_1661 % 6'h10; // @[util.scala 14:25:@225.4]
  assign _T_1662 = _GEN_22[4:0]; // @[util.scala 14:25:@225.4]
  assign _T_1663 = _T_1662 < _GEN_1139; // @[StoreQueue.scala 70:46:@226.4]
  assign initBits_7 = _T_1663 & io_bbStart; // @[StoreQueue.scala 70:64:@227.4]
  assign _T_1668 = 6'h18 - _GEN_1138; // @[util.scala 14:20:@229.4]
  assign _T_1669 = $unsigned(_T_1668); // @[util.scala 14:20:@230.4]
  assign _T_1670 = _T_1669[5:0]; // @[util.scala 14:20:@231.4]
  assign _GEN_23 = _T_1670 % 6'h10; // @[util.scala 14:25:@232.4]
  assign _T_1671 = _GEN_23[4:0]; // @[util.scala 14:25:@232.4]
  assign _T_1672 = _T_1671 < _GEN_1139; // @[StoreQueue.scala 70:46:@233.4]
  assign initBits_8 = _T_1672 & io_bbStart; // @[StoreQueue.scala 70:64:@234.4]
  assign _T_1677 = 6'h19 - _GEN_1138; // @[util.scala 14:20:@236.4]
  assign _T_1678 = $unsigned(_T_1677); // @[util.scala 14:20:@237.4]
  assign _T_1679 = _T_1678[5:0]; // @[util.scala 14:20:@238.4]
  assign _GEN_24 = _T_1679 % 6'h10; // @[util.scala 14:25:@239.4]
  assign _T_1680 = _GEN_24[4:0]; // @[util.scala 14:25:@239.4]
  assign _T_1681 = _T_1680 < _GEN_1139; // @[StoreQueue.scala 70:46:@240.4]
  assign initBits_9 = _T_1681 & io_bbStart; // @[StoreQueue.scala 70:64:@241.4]
  assign _T_1686 = 6'h1a - _GEN_1138; // @[util.scala 14:20:@243.4]
  assign _T_1687 = $unsigned(_T_1686); // @[util.scala 14:20:@244.4]
  assign _T_1688 = _T_1687[5:0]; // @[util.scala 14:20:@245.4]
  assign _GEN_25 = _T_1688 % 6'h10; // @[util.scala 14:25:@246.4]
  assign _T_1689 = _GEN_25[4:0]; // @[util.scala 14:25:@246.4]
  assign _T_1690 = _T_1689 < _GEN_1139; // @[StoreQueue.scala 70:46:@247.4]
  assign initBits_10 = _T_1690 & io_bbStart; // @[StoreQueue.scala 70:64:@248.4]
  assign _T_1695 = 6'h1b - _GEN_1138; // @[util.scala 14:20:@250.4]
  assign _T_1696 = $unsigned(_T_1695); // @[util.scala 14:20:@251.4]
  assign _T_1697 = _T_1696[5:0]; // @[util.scala 14:20:@252.4]
  assign _GEN_26 = _T_1697 % 6'h10; // @[util.scala 14:25:@253.4]
  assign _T_1698 = _GEN_26[4:0]; // @[util.scala 14:25:@253.4]
  assign _T_1699 = _T_1698 < _GEN_1139; // @[StoreQueue.scala 70:46:@254.4]
  assign initBits_11 = _T_1699 & io_bbStart; // @[StoreQueue.scala 70:64:@255.4]
  assign _T_1704 = 6'h1c - _GEN_1138; // @[util.scala 14:20:@257.4]
  assign _T_1705 = $unsigned(_T_1704); // @[util.scala 14:20:@258.4]
  assign _T_1706 = _T_1705[5:0]; // @[util.scala 14:20:@259.4]
  assign _GEN_27 = _T_1706 % 6'h10; // @[util.scala 14:25:@260.4]
  assign _T_1707 = _GEN_27[4:0]; // @[util.scala 14:25:@260.4]
  assign _T_1708 = _T_1707 < _GEN_1139; // @[StoreQueue.scala 70:46:@261.4]
  assign initBits_12 = _T_1708 & io_bbStart; // @[StoreQueue.scala 70:64:@262.4]
  assign _T_1713 = 6'h1d - _GEN_1138; // @[util.scala 14:20:@264.4]
  assign _T_1714 = $unsigned(_T_1713); // @[util.scala 14:20:@265.4]
  assign _T_1715 = _T_1714[5:0]; // @[util.scala 14:20:@266.4]
  assign _GEN_28 = _T_1715 % 6'h10; // @[util.scala 14:25:@267.4]
  assign _T_1716 = _GEN_28[4:0]; // @[util.scala 14:25:@267.4]
  assign _T_1717 = _T_1716 < _GEN_1139; // @[StoreQueue.scala 70:46:@268.4]
  assign initBits_13 = _T_1717 & io_bbStart; // @[StoreQueue.scala 70:64:@269.4]
  assign _T_1722 = 6'h1e - _GEN_1138; // @[util.scala 14:20:@271.4]
  assign _T_1723 = $unsigned(_T_1722); // @[util.scala 14:20:@272.4]
  assign _T_1724 = _T_1723[5:0]; // @[util.scala 14:20:@273.4]
  assign _GEN_29 = _T_1724 % 6'h10; // @[util.scala 14:25:@274.4]
  assign _T_1725 = _GEN_29[4:0]; // @[util.scala 14:25:@274.4]
  assign _T_1726 = _T_1725 < _GEN_1139; // @[StoreQueue.scala 70:46:@275.4]
  assign initBits_14 = _T_1726 & io_bbStart; // @[StoreQueue.scala 70:64:@276.4]
  assign _T_1731 = 6'h1f - _GEN_1138; // @[util.scala 14:20:@278.4]
  assign _T_1732 = $unsigned(_T_1731); // @[util.scala 14:20:@279.4]
  assign _T_1733 = _T_1732[5:0]; // @[util.scala 14:20:@280.4]
  assign _GEN_30 = _T_1733 % 6'h10; // @[util.scala 14:25:@281.4]
  assign _T_1734 = _GEN_30[4:0]; // @[util.scala 14:25:@281.4]
  assign _T_1735 = _T_1734 < _GEN_1139; // @[StoreQueue.scala 70:46:@282.4]
  assign initBits_15 = _T_1735 & io_bbStart; // @[StoreQueue.scala 70:64:@283.4]
  assign _T_1758 = allocatedEntries_0 | initBits_0; // @[StoreQueue.scala 72:78:@301.4]
  assign _T_1759 = allocatedEntries_1 | initBits_1; // @[StoreQueue.scala 72:78:@302.4]
  assign _T_1760 = allocatedEntries_2 | initBits_2; // @[StoreQueue.scala 72:78:@303.4]
  assign _T_1761 = allocatedEntries_3 | initBits_3; // @[StoreQueue.scala 72:78:@304.4]
  assign _T_1762 = allocatedEntries_4 | initBits_4; // @[StoreQueue.scala 72:78:@305.4]
  assign _T_1763 = allocatedEntries_5 | initBits_5; // @[StoreQueue.scala 72:78:@306.4]
  assign _T_1764 = allocatedEntries_6 | initBits_6; // @[StoreQueue.scala 72:78:@307.4]
  assign _T_1765 = allocatedEntries_7 | initBits_7; // @[StoreQueue.scala 72:78:@308.4]
  assign _T_1766 = allocatedEntries_8 | initBits_8; // @[StoreQueue.scala 72:78:@309.4]
  assign _T_1767 = allocatedEntries_9 | initBits_9; // @[StoreQueue.scala 72:78:@310.4]
  assign _T_1768 = allocatedEntries_10 | initBits_10; // @[StoreQueue.scala 72:78:@311.4]
  assign _T_1769 = allocatedEntries_11 | initBits_11; // @[StoreQueue.scala 72:78:@312.4]
  assign _T_1770 = allocatedEntries_12 | initBits_12; // @[StoreQueue.scala 72:78:@313.4]
  assign _T_1771 = allocatedEntries_13 | initBits_13; // @[StoreQueue.scala 72:78:@314.4]
  assign _T_1772 = allocatedEntries_14 | initBits_14; // @[StoreQueue.scala 72:78:@315.4]
  assign _T_1773 = allocatedEntries_15 | initBits_15; // @[StoreQueue.scala 72:78:@316.4]
  assign _T_1804 = _T_1599[3:0]; // @[:@356.6]
  assign _GEN_1 = 4'h1 == _T_1804 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_2 = 4'h2 == _T_1804 ? io_bbStoreOffsets_2 : _GEN_1; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_3 = 4'h3 == _T_1804 ? io_bbStoreOffsets_3 : _GEN_2; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_4 = 4'h4 == _T_1804 ? io_bbStoreOffsets_4 : _GEN_3; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_5 = 4'h5 == _T_1804 ? io_bbStoreOffsets_5 : _GEN_4; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_6 = 4'h6 == _T_1804 ? io_bbStoreOffsets_6 : _GEN_5; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_7 = 4'h7 == _T_1804 ? io_bbStoreOffsets_7 : _GEN_6; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_8 = 4'h8 == _T_1804 ? io_bbStoreOffsets_8 : _GEN_7; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_9 = 4'h9 == _T_1804 ? io_bbStoreOffsets_9 : _GEN_8; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_10 = 4'ha == _T_1804 ? io_bbStoreOffsets_10 : _GEN_9; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_11 = 4'hb == _T_1804 ? io_bbStoreOffsets_11 : _GEN_10; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_12 = 4'hc == _T_1804 ? io_bbStoreOffsets_12 : _GEN_11; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_13 = 4'hd == _T_1804 ? io_bbStoreOffsets_13 : _GEN_12; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_14 = 4'he == _T_1804 ? io_bbStoreOffsets_14 : _GEN_13; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_15 = 4'hf == _T_1804 ? io_bbStoreOffsets_15 : _GEN_14; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_32 = initBits_0 ? _GEN_15 : offsetQ_0; // @[StoreQueue.scala 75:25:@350.4]
  assign _GEN_33 = initBits_0 ? 1'h0 : portQ_0; // @[StoreQueue.scala 75:25:@350.4]
  assign _T_1822 = _T_1608[3:0]; // @[:@372.6]
  assign _GEN_35 = 4'h1 == _T_1822 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_36 = 4'h2 == _T_1822 ? io_bbStoreOffsets_2 : _GEN_35; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_37 = 4'h3 == _T_1822 ? io_bbStoreOffsets_3 : _GEN_36; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_38 = 4'h4 == _T_1822 ? io_bbStoreOffsets_4 : _GEN_37; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_39 = 4'h5 == _T_1822 ? io_bbStoreOffsets_5 : _GEN_38; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_40 = 4'h6 == _T_1822 ? io_bbStoreOffsets_6 : _GEN_39; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_41 = 4'h7 == _T_1822 ? io_bbStoreOffsets_7 : _GEN_40; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_42 = 4'h8 == _T_1822 ? io_bbStoreOffsets_8 : _GEN_41; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_43 = 4'h9 == _T_1822 ? io_bbStoreOffsets_9 : _GEN_42; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_44 = 4'ha == _T_1822 ? io_bbStoreOffsets_10 : _GEN_43; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_45 = 4'hb == _T_1822 ? io_bbStoreOffsets_11 : _GEN_44; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_46 = 4'hc == _T_1822 ? io_bbStoreOffsets_12 : _GEN_45; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_47 = 4'hd == _T_1822 ? io_bbStoreOffsets_13 : _GEN_46; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_48 = 4'he == _T_1822 ? io_bbStoreOffsets_14 : _GEN_47; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_49 = 4'hf == _T_1822 ? io_bbStoreOffsets_15 : _GEN_48; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_66 = initBits_1 ? _GEN_49 : offsetQ_1; // @[StoreQueue.scala 75:25:@366.4]
  assign _GEN_67 = initBits_1 ? 1'h0 : portQ_1; // @[StoreQueue.scala 75:25:@366.4]
  assign _T_1840 = _T_1617[3:0]; // @[:@388.6]
  assign _GEN_69 = 4'h1 == _T_1840 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_70 = 4'h2 == _T_1840 ? io_bbStoreOffsets_2 : _GEN_69; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_71 = 4'h3 == _T_1840 ? io_bbStoreOffsets_3 : _GEN_70; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_72 = 4'h4 == _T_1840 ? io_bbStoreOffsets_4 : _GEN_71; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_73 = 4'h5 == _T_1840 ? io_bbStoreOffsets_5 : _GEN_72; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_74 = 4'h6 == _T_1840 ? io_bbStoreOffsets_6 : _GEN_73; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_75 = 4'h7 == _T_1840 ? io_bbStoreOffsets_7 : _GEN_74; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_76 = 4'h8 == _T_1840 ? io_bbStoreOffsets_8 : _GEN_75; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_77 = 4'h9 == _T_1840 ? io_bbStoreOffsets_9 : _GEN_76; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_78 = 4'ha == _T_1840 ? io_bbStoreOffsets_10 : _GEN_77; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_79 = 4'hb == _T_1840 ? io_bbStoreOffsets_11 : _GEN_78; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_80 = 4'hc == _T_1840 ? io_bbStoreOffsets_12 : _GEN_79; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_81 = 4'hd == _T_1840 ? io_bbStoreOffsets_13 : _GEN_80; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_82 = 4'he == _T_1840 ? io_bbStoreOffsets_14 : _GEN_81; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_83 = 4'hf == _T_1840 ? io_bbStoreOffsets_15 : _GEN_82; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_100 = initBits_2 ? _GEN_83 : offsetQ_2; // @[StoreQueue.scala 75:25:@382.4]
  assign _GEN_101 = initBits_2 ? 1'h0 : portQ_2; // @[StoreQueue.scala 75:25:@382.4]
  assign _T_1858 = _T_1626[3:0]; // @[:@404.6]
  assign _GEN_103 = 4'h1 == _T_1858 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_104 = 4'h2 == _T_1858 ? io_bbStoreOffsets_2 : _GEN_103; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_105 = 4'h3 == _T_1858 ? io_bbStoreOffsets_3 : _GEN_104; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_106 = 4'h4 == _T_1858 ? io_bbStoreOffsets_4 : _GEN_105; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_107 = 4'h5 == _T_1858 ? io_bbStoreOffsets_5 : _GEN_106; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_108 = 4'h6 == _T_1858 ? io_bbStoreOffsets_6 : _GEN_107; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_109 = 4'h7 == _T_1858 ? io_bbStoreOffsets_7 : _GEN_108; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_110 = 4'h8 == _T_1858 ? io_bbStoreOffsets_8 : _GEN_109; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_111 = 4'h9 == _T_1858 ? io_bbStoreOffsets_9 : _GEN_110; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_112 = 4'ha == _T_1858 ? io_bbStoreOffsets_10 : _GEN_111; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_113 = 4'hb == _T_1858 ? io_bbStoreOffsets_11 : _GEN_112; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_114 = 4'hc == _T_1858 ? io_bbStoreOffsets_12 : _GEN_113; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_115 = 4'hd == _T_1858 ? io_bbStoreOffsets_13 : _GEN_114; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_116 = 4'he == _T_1858 ? io_bbStoreOffsets_14 : _GEN_115; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_117 = 4'hf == _T_1858 ? io_bbStoreOffsets_15 : _GEN_116; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_134 = initBits_3 ? _GEN_117 : offsetQ_3; // @[StoreQueue.scala 75:25:@398.4]
  assign _GEN_135 = initBits_3 ? 1'h0 : portQ_3; // @[StoreQueue.scala 75:25:@398.4]
  assign _T_1876 = _T_1635[3:0]; // @[:@420.6]
  assign _GEN_137 = 4'h1 == _T_1876 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_138 = 4'h2 == _T_1876 ? io_bbStoreOffsets_2 : _GEN_137; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_139 = 4'h3 == _T_1876 ? io_bbStoreOffsets_3 : _GEN_138; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_140 = 4'h4 == _T_1876 ? io_bbStoreOffsets_4 : _GEN_139; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_141 = 4'h5 == _T_1876 ? io_bbStoreOffsets_5 : _GEN_140; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_142 = 4'h6 == _T_1876 ? io_bbStoreOffsets_6 : _GEN_141; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_143 = 4'h7 == _T_1876 ? io_bbStoreOffsets_7 : _GEN_142; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_144 = 4'h8 == _T_1876 ? io_bbStoreOffsets_8 : _GEN_143; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_145 = 4'h9 == _T_1876 ? io_bbStoreOffsets_9 : _GEN_144; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_146 = 4'ha == _T_1876 ? io_bbStoreOffsets_10 : _GEN_145; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_147 = 4'hb == _T_1876 ? io_bbStoreOffsets_11 : _GEN_146; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_148 = 4'hc == _T_1876 ? io_bbStoreOffsets_12 : _GEN_147; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_149 = 4'hd == _T_1876 ? io_bbStoreOffsets_13 : _GEN_148; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_150 = 4'he == _T_1876 ? io_bbStoreOffsets_14 : _GEN_149; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_151 = 4'hf == _T_1876 ? io_bbStoreOffsets_15 : _GEN_150; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_168 = initBits_4 ? _GEN_151 : offsetQ_4; // @[StoreQueue.scala 75:25:@414.4]
  assign _GEN_169 = initBits_4 ? 1'h0 : portQ_4; // @[StoreQueue.scala 75:25:@414.4]
  assign _T_1894 = _T_1644[3:0]; // @[:@436.6]
  assign _GEN_171 = 4'h1 == _T_1894 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_172 = 4'h2 == _T_1894 ? io_bbStoreOffsets_2 : _GEN_171; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_173 = 4'h3 == _T_1894 ? io_bbStoreOffsets_3 : _GEN_172; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_174 = 4'h4 == _T_1894 ? io_bbStoreOffsets_4 : _GEN_173; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_175 = 4'h5 == _T_1894 ? io_bbStoreOffsets_5 : _GEN_174; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_176 = 4'h6 == _T_1894 ? io_bbStoreOffsets_6 : _GEN_175; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_177 = 4'h7 == _T_1894 ? io_bbStoreOffsets_7 : _GEN_176; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_178 = 4'h8 == _T_1894 ? io_bbStoreOffsets_8 : _GEN_177; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_179 = 4'h9 == _T_1894 ? io_bbStoreOffsets_9 : _GEN_178; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_180 = 4'ha == _T_1894 ? io_bbStoreOffsets_10 : _GEN_179; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_181 = 4'hb == _T_1894 ? io_bbStoreOffsets_11 : _GEN_180; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_182 = 4'hc == _T_1894 ? io_bbStoreOffsets_12 : _GEN_181; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_183 = 4'hd == _T_1894 ? io_bbStoreOffsets_13 : _GEN_182; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_184 = 4'he == _T_1894 ? io_bbStoreOffsets_14 : _GEN_183; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_185 = 4'hf == _T_1894 ? io_bbStoreOffsets_15 : _GEN_184; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_202 = initBits_5 ? _GEN_185 : offsetQ_5; // @[StoreQueue.scala 75:25:@430.4]
  assign _GEN_203 = initBits_5 ? 1'h0 : portQ_5; // @[StoreQueue.scala 75:25:@430.4]
  assign _T_1912 = _T_1653[3:0]; // @[:@452.6]
  assign _GEN_205 = 4'h1 == _T_1912 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_206 = 4'h2 == _T_1912 ? io_bbStoreOffsets_2 : _GEN_205; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_207 = 4'h3 == _T_1912 ? io_bbStoreOffsets_3 : _GEN_206; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_208 = 4'h4 == _T_1912 ? io_bbStoreOffsets_4 : _GEN_207; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_209 = 4'h5 == _T_1912 ? io_bbStoreOffsets_5 : _GEN_208; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_210 = 4'h6 == _T_1912 ? io_bbStoreOffsets_6 : _GEN_209; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_211 = 4'h7 == _T_1912 ? io_bbStoreOffsets_7 : _GEN_210; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_212 = 4'h8 == _T_1912 ? io_bbStoreOffsets_8 : _GEN_211; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_213 = 4'h9 == _T_1912 ? io_bbStoreOffsets_9 : _GEN_212; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_214 = 4'ha == _T_1912 ? io_bbStoreOffsets_10 : _GEN_213; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_215 = 4'hb == _T_1912 ? io_bbStoreOffsets_11 : _GEN_214; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_216 = 4'hc == _T_1912 ? io_bbStoreOffsets_12 : _GEN_215; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_217 = 4'hd == _T_1912 ? io_bbStoreOffsets_13 : _GEN_216; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_218 = 4'he == _T_1912 ? io_bbStoreOffsets_14 : _GEN_217; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_219 = 4'hf == _T_1912 ? io_bbStoreOffsets_15 : _GEN_218; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_236 = initBits_6 ? _GEN_219 : offsetQ_6; // @[StoreQueue.scala 75:25:@446.4]
  assign _GEN_237 = initBits_6 ? 1'h0 : portQ_6; // @[StoreQueue.scala 75:25:@446.4]
  assign _T_1930 = _T_1662[3:0]; // @[:@468.6]
  assign _GEN_239 = 4'h1 == _T_1930 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_240 = 4'h2 == _T_1930 ? io_bbStoreOffsets_2 : _GEN_239; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_241 = 4'h3 == _T_1930 ? io_bbStoreOffsets_3 : _GEN_240; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_242 = 4'h4 == _T_1930 ? io_bbStoreOffsets_4 : _GEN_241; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_243 = 4'h5 == _T_1930 ? io_bbStoreOffsets_5 : _GEN_242; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_244 = 4'h6 == _T_1930 ? io_bbStoreOffsets_6 : _GEN_243; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_245 = 4'h7 == _T_1930 ? io_bbStoreOffsets_7 : _GEN_244; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_246 = 4'h8 == _T_1930 ? io_bbStoreOffsets_8 : _GEN_245; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_247 = 4'h9 == _T_1930 ? io_bbStoreOffsets_9 : _GEN_246; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_248 = 4'ha == _T_1930 ? io_bbStoreOffsets_10 : _GEN_247; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_249 = 4'hb == _T_1930 ? io_bbStoreOffsets_11 : _GEN_248; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_250 = 4'hc == _T_1930 ? io_bbStoreOffsets_12 : _GEN_249; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_251 = 4'hd == _T_1930 ? io_bbStoreOffsets_13 : _GEN_250; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_252 = 4'he == _T_1930 ? io_bbStoreOffsets_14 : _GEN_251; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_253 = 4'hf == _T_1930 ? io_bbStoreOffsets_15 : _GEN_252; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_270 = initBits_7 ? _GEN_253 : offsetQ_7; // @[StoreQueue.scala 75:25:@462.4]
  assign _GEN_271 = initBits_7 ? 1'h0 : portQ_7; // @[StoreQueue.scala 75:25:@462.4]
  assign _T_1948 = _T_1671[3:0]; // @[:@484.6]
  assign _GEN_273 = 4'h1 == _T_1948 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_274 = 4'h2 == _T_1948 ? io_bbStoreOffsets_2 : _GEN_273; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_275 = 4'h3 == _T_1948 ? io_bbStoreOffsets_3 : _GEN_274; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_276 = 4'h4 == _T_1948 ? io_bbStoreOffsets_4 : _GEN_275; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_277 = 4'h5 == _T_1948 ? io_bbStoreOffsets_5 : _GEN_276; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_278 = 4'h6 == _T_1948 ? io_bbStoreOffsets_6 : _GEN_277; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_279 = 4'h7 == _T_1948 ? io_bbStoreOffsets_7 : _GEN_278; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_280 = 4'h8 == _T_1948 ? io_bbStoreOffsets_8 : _GEN_279; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_281 = 4'h9 == _T_1948 ? io_bbStoreOffsets_9 : _GEN_280; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_282 = 4'ha == _T_1948 ? io_bbStoreOffsets_10 : _GEN_281; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_283 = 4'hb == _T_1948 ? io_bbStoreOffsets_11 : _GEN_282; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_284 = 4'hc == _T_1948 ? io_bbStoreOffsets_12 : _GEN_283; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_285 = 4'hd == _T_1948 ? io_bbStoreOffsets_13 : _GEN_284; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_286 = 4'he == _T_1948 ? io_bbStoreOffsets_14 : _GEN_285; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_287 = 4'hf == _T_1948 ? io_bbStoreOffsets_15 : _GEN_286; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_304 = initBits_8 ? _GEN_287 : offsetQ_8; // @[StoreQueue.scala 75:25:@478.4]
  assign _GEN_305 = initBits_8 ? 1'h0 : portQ_8; // @[StoreQueue.scala 75:25:@478.4]
  assign _T_1966 = _T_1680[3:0]; // @[:@500.6]
  assign _GEN_307 = 4'h1 == _T_1966 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_308 = 4'h2 == _T_1966 ? io_bbStoreOffsets_2 : _GEN_307; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_309 = 4'h3 == _T_1966 ? io_bbStoreOffsets_3 : _GEN_308; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_310 = 4'h4 == _T_1966 ? io_bbStoreOffsets_4 : _GEN_309; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_311 = 4'h5 == _T_1966 ? io_bbStoreOffsets_5 : _GEN_310; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_312 = 4'h6 == _T_1966 ? io_bbStoreOffsets_6 : _GEN_311; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_313 = 4'h7 == _T_1966 ? io_bbStoreOffsets_7 : _GEN_312; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_314 = 4'h8 == _T_1966 ? io_bbStoreOffsets_8 : _GEN_313; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_315 = 4'h9 == _T_1966 ? io_bbStoreOffsets_9 : _GEN_314; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_316 = 4'ha == _T_1966 ? io_bbStoreOffsets_10 : _GEN_315; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_317 = 4'hb == _T_1966 ? io_bbStoreOffsets_11 : _GEN_316; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_318 = 4'hc == _T_1966 ? io_bbStoreOffsets_12 : _GEN_317; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_319 = 4'hd == _T_1966 ? io_bbStoreOffsets_13 : _GEN_318; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_320 = 4'he == _T_1966 ? io_bbStoreOffsets_14 : _GEN_319; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_321 = 4'hf == _T_1966 ? io_bbStoreOffsets_15 : _GEN_320; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_338 = initBits_9 ? _GEN_321 : offsetQ_9; // @[StoreQueue.scala 75:25:@494.4]
  assign _GEN_339 = initBits_9 ? 1'h0 : portQ_9; // @[StoreQueue.scala 75:25:@494.4]
  assign _T_1984 = _T_1689[3:0]; // @[:@516.6]
  assign _GEN_341 = 4'h1 == _T_1984 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_342 = 4'h2 == _T_1984 ? io_bbStoreOffsets_2 : _GEN_341; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_343 = 4'h3 == _T_1984 ? io_bbStoreOffsets_3 : _GEN_342; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_344 = 4'h4 == _T_1984 ? io_bbStoreOffsets_4 : _GEN_343; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_345 = 4'h5 == _T_1984 ? io_bbStoreOffsets_5 : _GEN_344; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_346 = 4'h6 == _T_1984 ? io_bbStoreOffsets_6 : _GEN_345; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_347 = 4'h7 == _T_1984 ? io_bbStoreOffsets_7 : _GEN_346; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_348 = 4'h8 == _T_1984 ? io_bbStoreOffsets_8 : _GEN_347; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_349 = 4'h9 == _T_1984 ? io_bbStoreOffsets_9 : _GEN_348; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_350 = 4'ha == _T_1984 ? io_bbStoreOffsets_10 : _GEN_349; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_351 = 4'hb == _T_1984 ? io_bbStoreOffsets_11 : _GEN_350; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_352 = 4'hc == _T_1984 ? io_bbStoreOffsets_12 : _GEN_351; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_353 = 4'hd == _T_1984 ? io_bbStoreOffsets_13 : _GEN_352; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_354 = 4'he == _T_1984 ? io_bbStoreOffsets_14 : _GEN_353; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_355 = 4'hf == _T_1984 ? io_bbStoreOffsets_15 : _GEN_354; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_372 = initBits_10 ? _GEN_355 : offsetQ_10; // @[StoreQueue.scala 75:25:@510.4]
  assign _GEN_373 = initBits_10 ? 1'h0 : portQ_10; // @[StoreQueue.scala 75:25:@510.4]
  assign _T_2002 = _T_1698[3:0]; // @[:@532.6]
  assign _GEN_375 = 4'h1 == _T_2002 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_376 = 4'h2 == _T_2002 ? io_bbStoreOffsets_2 : _GEN_375; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_377 = 4'h3 == _T_2002 ? io_bbStoreOffsets_3 : _GEN_376; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_378 = 4'h4 == _T_2002 ? io_bbStoreOffsets_4 : _GEN_377; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_379 = 4'h5 == _T_2002 ? io_bbStoreOffsets_5 : _GEN_378; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_380 = 4'h6 == _T_2002 ? io_bbStoreOffsets_6 : _GEN_379; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_381 = 4'h7 == _T_2002 ? io_bbStoreOffsets_7 : _GEN_380; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_382 = 4'h8 == _T_2002 ? io_bbStoreOffsets_8 : _GEN_381; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_383 = 4'h9 == _T_2002 ? io_bbStoreOffsets_9 : _GEN_382; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_384 = 4'ha == _T_2002 ? io_bbStoreOffsets_10 : _GEN_383; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_385 = 4'hb == _T_2002 ? io_bbStoreOffsets_11 : _GEN_384; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_386 = 4'hc == _T_2002 ? io_bbStoreOffsets_12 : _GEN_385; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_387 = 4'hd == _T_2002 ? io_bbStoreOffsets_13 : _GEN_386; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_388 = 4'he == _T_2002 ? io_bbStoreOffsets_14 : _GEN_387; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_389 = 4'hf == _T_2002 ? io_bbStoreOffsets_15 : _GEN_388; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_406 = initBits_11 ? _GEN_389 : offsetQ_11; // @[StoreQueue.scala 75:25:@526.4]
  assign _GEN_407 = initBits_11 ? 1'h0 : portQ_11; // @[StoreQueue.scala 75:25:@526.4]
  assign _T_2020 = _T_1707[3:0]; // @[:@548.6]
  assign _GEN_409 = 4'h1 == _T_2020 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_410 = 4'h2 == _T_2020 ? io_bbStoreOffsets_2 : _GEN_409; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_411 = 4'h3 == _T_2020 ? io_bbStoreOffsets_3 : _GEN_410; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_412 = 4'h4 == _T_2020 ? io_bbStoreOffsets_4 : _GEN_411; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_413 = 4'h5 == _T_2020 ? io_bbStoreOffsets_5 : _GEN_412; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_414 = 4'h6 == _T_2020 ? io_bbStoreOffsets_6 : _GEN_413; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_415 = 4'h7 == _T_2020 ? io_bbStoreOffsets_7 : _GEN_414; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_416 = 4'h8 == _T_2020 ? io_bbStoreOffsets_8 : _GEN_415; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_417 = 4'h9 == _T_2020 ? io_bbStoreOffsets_9 : _GEN_416; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_418 = 4'ha == _T_2020 ? io_bbStoreOffsets_10 : _GEN_417; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_419 = 4'hb == _T_2020 ? io_bbStoreOffsets_11 : _GEN_418; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_420 = 4'hc == _T_2020 ? io_bbStoreOffsets_12 : _GEN_419; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_421 = 4'hd == _T_2020 ? io_bbStoreOffsets_13 : _GEN_420; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_422 = 4'he == _T_2020 ? io_bbStoreOffsets_14 : _GEN_421; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_423 = 4'hf == _T_2020 ? io_bbStoreOffsets_15 : _GEN_422; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_440 = initBits_12 ? _GEN_423 : offsetQ_12; // @[StoreQueue.scala 75:25:@542.4]
  assign _GEN_441 = initBits_12 ? 1'h0 : portQ_12; // @[StoreQueue.scala 75:25:@542.4]
  assign _T_2038 = _T_1716[3:0]; // @[:@564.6]
  assign _GEN_443 = 4'h1 == _T_2038 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_444 = 4'h2 == _T_2038 ? io_bbStoreOffsets_2 : _GEN_443; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_445 = 4'h3 == _T_2038 ? io_bbStoreOffsets_3 : _GEN_444; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_446 = 4'h4 == _T_2038 ? io_bbStoreOffsets_4 : _GEN_445; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_447 = 4'h5 == _T_2038 ? io_bbStoreOffsets_5 : _GEN_446; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_448 = 4'h6 == _T_2038 ? io_bbStoreOffsets_6 : _GEN_447; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_449 = 4'h7 == _T_2038 ? io_bbStoreOffsets_7 : _GEN_448; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_450 = 4'h8 == _T_2038 ? io_bbStoreOffsets_8 : _GEN_449; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_451 = 4'h9 == _T_2038 ? io_bbStoreOffsets_9 : _GEN_450; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_452 = 4'ha == _T_2038 ? io_bbStoreOffsets_10 : _GEN_451; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_453 = 4'hb == _T_2038 ? io_bbStoreOffsets_11 : _GEN_452; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_454 = 4'hc == _T_2038 ? io_bbStoreOffsets_12 : _GEN_453; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_455 = 4'hd == _T_2038 ? io_bbStoreOffsets_13 : _GEN_454; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_456 = 4'he == _T_2038 ? io_bbStoreOffsets_14 : _GEN_455; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_457 = 4'hf == _T_2038 ? io_bbStoreOffsets_15 : _GEN_456; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_474 = initBits_13 ? _GEN_457 : offsetQ_13; // @[StoreQueue.scala 75:25:@558.4]
  assign _GEN_475 = initBits_13 ? 1'h0 : portQ_13; // @[StoreQueue.scala 75:25:@558.4]
  assign _T_2056 = _T_1725[3:0]; // @[:@580.6]
  assign _GEN_477 = 4'h1 == _T_2056 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_478 = 4'h2 == _T_2056 ? io_bbStoreOffsets_2 : _GEN_477; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_479 = 4'h3 == _T_2056 ? io_bbStoreOffsets_3 : _GEN_478; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_480 = 4'h4 == _T_2056 ? io_bbStoreOffsets_4 : _GEN_479; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_481 = 4'h5 == _T_2056 ? io_bbStoreOffsets_5 : _GEN_480; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_482 = 4'h6 == _T_2056 ? io_bbStoreOffsets_6 : _GEN_481; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_483 = 4'h7 == _T_2056 ? io_bbStoreOffsets_7 : _GEN_482; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_484 = 4'h8 == _T_2056 ? io_bbStoreOffsets_8 : _GEN_483; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_485 = 4'h9 == _T_2056 ? io_bbStoreOffsets_9 : _GEN_484; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_486 = 4'ha == _T_2056 ? io_bbStoreOffsets_10 : _GEN_485; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_487 = 4'hb == _T_2056 ? io_bbStoreOffsets_11 : _GEN_486; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_488 = 4'hc == _T_2056 ? io_bbStoreOffsets_12 : _GEN_487; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_489 = 4'hd == _T_2056 ? io_bbStoreOffsets_13 : _GEN_488; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_490 = 4'he == _T_2056 ? io_bbStoreOffsets_14 : _GEN_489; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_491 = 4'hf == _T_2056 ? io_bbStoreOffsets_15 : _GEN_490; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_508 = initBits_14 ? _GEN_491 : offsetQ_14; // @[StoreQueue.scala 75:25:@574.4]
  assign _GEN_509 = initBits_14 ? 1'h0 : portQ_14; // @[StoreQueue.scala 75:25:@574.4]
  assign _T_2074 = _T_1734[3:0]; // @[:@596.6]
  assign _GEN_511 = 4'h1 == _T_2074 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_512 = 4'h2 == _T_2074 ? io_bbStoreOffsets_2 : _GEN_511; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_513 = 4'h3 == _T_2074 ? io_bbStoreOffsets_3 : _GEN_512; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_514 = 4'h4 == _T_2074 ? io_bbStoreOffsets_4 : _GEN_513; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_515 = 4'h5 == _T_2074 ? io_bbStoreOffsets_5 : _GEN_514; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_516 = 4'h6 == _T_2074 ? io_bbStoreOffsets_6 : _GEN_515; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_517 = 4'h7 == _T_2074 ? io_bbStoreOffsets_7 : _GEN_516; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_518 = 4'h8 == _T_2074 ? io_bbStoreOffsets_8 : _GEN_517; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_519 = 4'h9 == _T_2074 ? io_bbStoreOffsets_9 : _GEN_518; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_520 = 4'ha == _T_2074 ? io_bbStoreOffsets_10 : _GEN_519; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_521 = 4'hb == _T_2074 ? io_bbStoreOffsets_11 : _GEN_520; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_522 = 4'hc == _T_2074 ? io_bbStoreOffsets_12 : _GEN_521; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_523 = 4'hd == _T_2074 ? io_bbStoreOffsets_13 : _GEN_522; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_524 = 4'he == _T_2074 ? io_bbStoreOffsets_14 : _GEN_523; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_525 = 4'hf == _T_2074 ? io_bbStoreOffsets_15 : _GEN_524; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_542 = initBits_15 ? _GEN_525 : offsetQ_15; // @[StoreQueue.scala 75:25:@590.4]
  assign _GEN_543 = initBits_15 ? 1'h0 : portQ_15; // @[StoreQueue.scala 75:25:@590.4]
  assign _T_2096 = _GEN_15 + 4'h1; // @[util.scala 10:8:@615.6]
  assign _GEN_31 = _T_2096 % 5'h10; // @[util.scala 10:14:@616.6]
  assign _T_2097 = _GEN_31[4:0]; // @[util.scala 10:14:@616.6]
  assign _GEN_1203 = {{1'd0}, io_loadTail}; // @[StoreQueue.scala 96:56:@617.6]
  assign _T_2098 = _T_2097 == _GEN_1203; // @[StoreQueue.scala 96:56:@617.6]
  assign _T_2099 = io_loadEmpty & _T_2098; // @[StoreQueue.scala 95:50:@618.6]
  assign _T_2101 = _T_2099 == 1'h0; // @[StoreQueue.scala 95:35:@619.6]
  assign _T_2103 = previousLoadHead <= offsetQ_0; // @[StoreQueue.scala 100:35:@627.8]
  assign _T_2104 = offsetQ_0 < io_loadHead; // @[StoreQueue.scala 100:87:@628.8]
  assign _T_2105 = _T_2103 & _T_2104; // @[StoreQueue.scala 100:61:@629.8]
  assign _T_2107 = previousLoadHead > io_loadHead; // @[StoreQueue.scala 102:35:@634.10]
  assign _T_2108 = io_loadHead <= offsetQ_0; // @[StoreQueue.scala 103:23:@635.10]
  assign _T_2109 = offsetQ_0 < previousLoadHead; // @[StoreQueue.scala 103:75:@636.10]
  assign _T_2110 = _T_2108 & _T_2109; // @[StoreQueue.scala 103:49:@637.10]
  assign _T_2112 = _T_2110 == 1'h0; // @[StoreQueue.scala 103:9:@638.10]
  assign _T_2113 = _T_2107 & _T_2112; // @[StoreQueue.scala 102:49:@639.10]
  assign _GEN_560 = _T_2113 ? 1'h0 : checkBits_0; // @[StoreQueue.scala 103:96:@640.10]
  assign _GEN_561 = _T_2105 ? 1'h0 : _GEN_560; // @[StoreQueue.scala 100:102:@630.8]
  assign _GEN_562 = io_loadEmpty ? 1'h0 : _GEN_561; // @[StoreQueue.scala 98:26:@623.6]
  assign _GEN_563 = initBits_0 ? _T_2101 : _GEN_562; // @[StoreQueue.scala 94:35:@608.4]
  assign _T_2126 = _GEN_49 + 4'h1; // @[util.scala 10:8:@651.6]
  assign _GEN_34 = _T_2126 % 5'h10; // @[util.scala 10:14:@652.6]
  assign _T_2127 = _GEN_34[4:0]; // @[util.scala 10:14:@652.6]
  assign _T_2128 = _T_2127 == _GEN_1203; // @[StoreQueue.scala 96:56:@653.6]
  assign _T_2129 = io_loadEmpty & _T_2128; // @[StoreQueue.scala 95:50:@654.6]
  assign _T_2131 = _T_2129 == 1'h0; // @[StoreQueue.scala 95:35:@655.6]
  assign _T_2133 = previousLoadHead <= offsetQ_1; // @[StoreQueue.scala 100:35:@663.8]
  assign _T_2134 = offsetQ_1 < io_loadHead; // @[StoreQueue.scala 100:87:@664.8]
  assign _T_2135 = _T_2133 & _T_2134; // @[StoreQueue.scala 100:61:@665.8]
  assign _T_2138 = io_loadHead <= offsetQ_1; // @[StoreQueue.scala 103:23:@671.10]
  assign _T_2139 = offsetQ_1 < previousLoadHead; // @[StoreQueue.scala 103:75:@672.10]
  assign _T_2140 = _T_2138 & _T_2139; // @[StoreQueue.scala 103:49:@673.10]
  assign _T_2142 = _T_2140 == 1'h0; // @[StoreQueue.scala 103:9:@674.10]
  assign _T_2143 = _T_2107 & _T_2142; // @[StoreQueue.scala 102:49:@675.10]
  assign _GEN_580 = _T_2143 ? 1'h0 : checkBits_1; // @[StoreQueue.scala 103:96:@676.10]
  assign _GEN_581 = _T_2135 ? 1'h0 : _GEN_580; // @[StoreQueue.scala 100:102:@666.8]
  assign _GEN_582 = io_loadEmpty ? 1'h0 : _GEN_581; // @[StoreQueue.scala 98:26:@659.6]
  assign _GEN_583 = initBits_1 ? _T_2131 : _GEN_582; // @[StoreQueue.scala 94:35:@644.4]
  assign _T_2156 = _GEN_83 + 4'h1; // @[util.scala 10:8:@687.6]
  assign _GEN_50 = _T_2156 % 5'h10; // @[util.scala 10:14:@688.6]
  assign _T_2157 = _GEN_50[4:0]; // @[util.scala 10:14:@688.6]
  assign _T_2158 = _T_2157 == _GEN_1203; // @[StoreQueue.scala 96:56:@689.6]
  assign _T_2159 = io_loadEmpty & _T_2158; // @[StoreQueue.scala 95:50:@690.6]
  assign _T_2161 = _T_2159 == 1'h0; // @[StoreQueue.scala 95:35:@691.6]
  assign _T_2163 = previousLoadHead <= offsetQ_2; // @[StoreQueue.scala 100:35:@699.8]
  assign _T_2164 = offsetQ_2 < io_loadHead; // @[StoreQueue.scala 100:87:@700.8]
  assign _T_2165 = _T_2163 & _T_2164; // @[StoreQueue.scala 100:61:@701.8]
  assign _T_2168 = io_loadHead <= offsetQ_2; // @[StoreQueue.scala 103:23:@707.10]
  assign _T_2169 = offsetQ_2 < previousLoadHead; // @[StoreQueue.scala 103:75:@708.10]
  assign _T_2170 = _T_2168 & _T_2169; // @[StoreQueue.scala 103:49:@709.10]
  assign _T_2172 = _T_2170 == 1'h0; // @[StoreQueue.scala 103:9:@710.10]
  assign _T_2173 = _T_2107 & _T_2172; // @[StoreQueue.scala 102:49:@711.10]
  assign _GEN_600 = _T_2173 ? 1'h0 : checkBits_2; // @[StoreQueue.scala 103:96:@712.10]
  assign _GEN_601 = _T_2165 ? 1'h0 : _GEN_600; // @[StoreQueue.scala 100:102:@702.8]
  assign _GEN_602 = io_loadEmpty ? 1'h0 : _GEN_601; // @[StoreQueue.scala 98:26:@695.6]
  assign _GEN_603 = initBits_2 ? _T_2161 : _GEN_602; // @[StoreQueue.scala 94:35:@680.4]
  assign _T_2186 = _GEN_117 + 4'h1; // @[util.scala 10:8:@723.6]
  assign _GEN_51 = _T_2186 % 5'h10; // @[util.scala 10:14:@724.6]
  assign _T_2187 = _GEN_51[4:0]; // @[util.scala 10:14:@724.6]
  assign _T_2188 = _T_2187 == _GEN_1203; // @[StoreQueue.scala 96:56:@725.6]
  assign _T_2189 = io_loadEmpty & _T_2188; // @[StoreQueue.scala 95:50:@726.6]
  assign _T_2191 = _T_2189 == 1'h0; // @[StoreQueue.scala 95:35:@727.6]
  assign _T_2193 = previousLoadHead <= offsetQ_3; // @[StoreQueue.scala 100:35:@735.8]
  assign _T_2194 = offsetQ_3 < io_loadHead; // @[StoreQueue.scala 100:87:@736.8]
  assign _T_2195 = _T_2193 & _T_2194; // @[StoreQueue.scala 100:61:@737.8]
  assign _T_2198 = io_loadHead <= offsetQ_3; // @[StoreQueue.scala 103:23:@743.10]
  assign _T_2199 = offsetQ_3 < previousLoadHead; // @[StoreQueue.scala 103:75:@744.10]
  assign _T_2200 = _T_2198 & _T_2199; // @[StoreQueue.scala 103:49:@745.10]
  assign _T_2202 = _T_2200 == 1'h0; // @[StoreQueue.scala 103:9:@746.10]
  assign _T_2203 = _T_2107 & _T_2202; // @[StoreQueue.scala 102:49:@747.10]
  assign _GEN_620 = _T_2203 ? 1'h0 : checkBits_3; // @[StoreQueue.scala 103:96:@748.10]
  assign _GEN_621 = _T_2195 ? 1'h0 : _GEN_620; // @[StoreQueue.scala 100:102:@738.8]
  assign _GEN_622 = io_loadEmpty ? 1'h0 : _GEN_621; // @[StoreQueue.scala 98:26:@731.6]
  assign _GEN_623 = initBits_3 ? _T_2191 : _GEN_622; // @[StoreQueue.scala 94:35:@716.4]
  assign _T_2216 = _GEN_151 + 4'h1; // @[util.scala 10:8:@759.6]
  assign _GEN_52 = _T_2216 % 5'h10; // @[util.scala 10:14:@760.6]
  assign _T_2217 = _GEN_52[4:0]; // @[util.scala 10:14:@760.6]
  assign _T_2218 = _T_2217 == _GEN_1203; // @[StoreQueue.scala 96:56:@761.6]
  assign _T_2219 = io_loadEmpty & _T_2218; // @[StoreQueue.scala 95:50:@762.6]
  assign _T_2221 = _T_2219 == 1'h0; // @[StoreQueue.scala 95:35:@763.6]
  assign _T_2223 = previousLoadHead <= offsetQ_4; // @[StoreQueue.scala 100:35:@771.8]
  assign _T_2224 = offsetQ_4 < io_loadHead; // @[StoreQueue.scala 100:87:@772.8]
  assign _T_2225 = _T_2223 & _T_2224; // @[StoreQueue.scala 100:61:@773.8]
  assign _T_2228 = io_loadHead <= offsetQ_4; // @[StoreQueue.scala 103:23:@779.10]
  assign _T_2229 = offsetQ_4 < previousLoadHead; // @[StoreQueue.scala 103:75:@780.10]
  assign _T_2230 = _T_2228 & _T_2229; // @[StoreQueue.scala 103:49:@781.10]
  assign _T_2232 = _T_2230 == 1'h0; // @[StoreQueue.scala 103:9:@782.10]
  assign _T_2233 = _T_2107 & _T_2232; // @[StoreQueue.scala 102:49:@783.10]
  assign _GEN_640 = _T_2233 ? 1'h0 : checkBits_4; // @[StoreQueue.scala 103:96:@784.10]
  assign _GEN_641 = _T_2225 ? 1'h0 : _GEN_640; // @[StoreQueue.scala 100:102:@774.8]
  assign _GEN_642 = io_loadEmpty ? 1'h0 : _GEN_641; // @[StoreQueue.scala 98:26:@767.6]
  assign _GEN_643 = initBits_4 ? _T_2221 : _GEN_642; // @[StoreQueue.scala 94:35:@752.4]
  assign _T_2246 = _GEN_185 + 4'h1; // @[util.scala 10:8:@795.6]
  assign _GEN_53 = _T_2246 % 5'h10; // @[util.scala 10:14:@796.6]
  assign _T_2247 = _GEN_53[4:0]; // @[util.scala 10:14:@796.6]
  assign _T_2248 = _T_2247 == _GEN_1203; // @[StoreQueue.scala 96:56:@797.6]
  assign _T_2249 = io_loadEmpty & _T_2248; // @[StoreQueue.scala 95:50:@798.6]
  assign _T_2251 = _T_2249 == 1'h0; // @[StoreQueue.scala 95:35:@799.6]
  assign _T_2253 = previousLoadHead <= offsetQ_5; // @[StoreQueue.scala 100:35:@807.8]
  assign _T_2254 = offsetQ_5 < io_loadHead; // @[StoreQueue.scala 100:87:@808.8]
  assign _T_2255 = _T_2253 & _T_2254; // @[StoreQueue.scala 100:61:@809.8]
  assign _T_2258 = io_loadHead <= offsetQ_5; // @[StoreQueue.scala 103:23:@815.10]
  assign _T_2259 = offsetQ_5 < previousLoadHead; // @[StoreQueue.scala 103:75:@816.10]
  assign _T_2260 = _T_2258 & _T_2259; // @[StoreQueue.scala 103:49:@817.10]
  assign _T_2262 = _T_2260 == 1'h0; // @[StoreQueue.scala 103:9:@818.10]
  assign _T_2263 = _T_2107 & _T_2262; // @[StoreQueue.scala 102:49:@819.10]
  assign _GEN_660 = _T_2263 ? 1'h0 : checkBits_5; // @[StoreQueue.scala 103:96:@820.10]
  assign _GEN_661 = _T_2255 ? 1'h0 : _GEN_660; // @[StoreQueue.scala 100:102:@810.8]
  assign _GEN_662 = io_loadEmpty ? 1'h0 : _GEN_661; // @[StoreQueue.scala 98:26:@803.6]
  assign _GEN_663 = initBits_5 ? _T_2251 : _GEN_662; // @[StoreQueue.scala 94:35:@788.4]
  assign _T_2276 = _GEN_219 + 4'h1; // @[util.scala 10:8:@831.6]
  assign _GEN_54 = _T_2276 % 5'h10; // @[util.scala 10:14:@832.6]
  assign _T_2277 = _GEN_54[4:0]; // @[util.scala 10:14:@832.6]
  assign _T_2278 = _T_2277 == _GEN_1203; // @[StoreQueue.scala 96:56:@833.6]
  assign _T_2279 = io_loadEmpty & _T_2278; // @[StoreQueue.scala 95:50:@834.6]
  assign _T_2281 = _T_2279 == 1'h0; // @[StoreQueue.scala 95:35:@835.6]
  assign _T_2283 = previousLoadHead <= offsetQ_6; // @[StoreQueue.scala 100:35:@843.8]
  assign _T_2284 = offsetQ_6 < io_loadHead; // @[StoreQueue.scala 100:87:@844.8]
  assign _T_2285 = _T_2283 & _T_2284; // @[StoreQueue.scala 100:61:@845.8]
  assign _T_2288 = io_loadHead <= offsetQ_6; // @[StoreQueue.scala 103:23:@851.10]
  assign _T_2289 = offsetQ_6 < previousLoadHead; // @[StoreQueue.scala 103:75:@852.10]
  assign _T_2290 = _T_2288 & _T_2289; // @[StoreQueue.scala 103:49:@853.10]
  assign _T_2292 = _T_2290 == 1'h0; // @[StoreQueue.scala 103:9:@854.10]
  assign _T_2293 = _T_2107 & _T_2292; // @[StoreQueue.scala 102:49:@855.10]
  assign _GEN_680 = _T_2293 ? 1'h0 : checkBits_6; // @[StoreQueue.scala 103:96:@856.10]
  assign _GEN_681 = _T_2285 ? 1'h0 : _GEN_680; // @[StoreQueue.scala 100:102:@846.8]
  assign _GEN_682 = io_loadEmpty ? 1'h0 : _GEN_681; // @[StoreQueue.scala 98:26:@839.6]
  assign _GEN_683 = initBits_6 ? _T_2281 : _GEN_682; // @[StoreQueue.scala 94:35:@824.4]
  assign _T_2306 = _GEN_253 + 4'h1; // @[util.scala 10:8:@867.6]
  assign _GEN_55 = _T_2306 % 5'h10; // @[util.scala 10:14:@868.6]
  assign _T_2307 = _GEN_55[4:0]; // @[util.scala 10:14:@868.6]
  assign _T_2308 = _T_2307 == _GEN_1203; // @[StoreQueue.scala 96:56:@869.6]
  assign _T_2309 = io_loadEmpty & _T_2308; // @[StoreQueue.scala 95:50:@870.6]
  assign _T_2311 = _T_2309 == 1'h0; // @[StoreQueue.scala 95:35:@871.6]
  assign _T_2313 = previousLoadHead <= offsetQ_7; // @[StoreQueue.scala 100:35:@879.8]
  assign _T_2314 = offsetQ_7 < io_loadHead; // @[StoreQueue.scala 100:87:@880.8]
  assign _T_2315 = _T_2313 & _T_2314; // @[StoreQueue.scala 100:61:@881.8]
  assign _T_2318 = io_loadHead <= offsetQ_7; // @[StoreQueue.scala 103:23:@887.10]
  assign _T_2319 = offsetQ_7 < previousLoadHead; // @[StoreQueue.scala 103:75:@888.10]
  assign _T_2320 = _T_2318 & _T_2319; // @[StoreQueue.scala 103:49:@889.10]
  assign _T_2322 = _T_2320 == 1'h0; // @[StoreQueue.scala 103:9:@890.10]
  assign _T_2323 = _T_2107 & _T_2322; // @[StoreQueue.scala 102:49:@891.10]
  assign _GEN_700 = _T_2323 ? 1'h0 : checkBits_7; // @[StoreQueue.scala 103:96:@892.10]
  assign _GEN_701 = _T_2315 ? 1'h0 : _GEN_700; // @[StoreQueue.scala 100:102:@882.8]
  assign _GEN_702 = io_loadEmpty ? 1'h0 : _GEN_701; // @[StoreQueue.scala 98:26:@875.6]
  assign _GEN_703 = initBits_7 ? _T_2311 : _GEN_702; // @[StoreQueue.scala 94:35:@860.4]
  assign _T_2336 = _GEN_287 + 4'h1; // @[util.scala 10:8:@903.6]
  assign _GEN_56 = _T_2336 % 5'h10; // @[util.scala 10:14:@904.6]
  assign _T_2337 = _GEN_56[4:0]; // @[util.scala 10:14:@904.6]
  assign _T_2338 = _T_2337 == _GEN_1203; // @[StoreQueue.scala 96:56:@905.6]
  assign _T_2339 = io_loadEmpty & _T_2338; // @[StoreQueue.scala 95:50:@906.6]
  assign _T_2341 = _T_2339 == 1'h0; // @[StoreQueue.scala 95:35:@907.6]
  assign _T_2343 = previousLoadHead <= offsetQ_8; // @[StoreQueue.scala 100:35:@915.8]
  assign _T_2344 = offsetQ_8 < io_loadHead; // @[StoreQueue.scala 100:87:@916.8]
  assign _T_2345 = _T_2343 & _T_2344; // @[StoreQueue.scala 100:61:@917.8]
  assign _T_2348 = io_loadHead <= offsetQ_8; // @[StoreQueue.scala 103:23:@923.10]
  assign _T_2349 = offsetQ_8 < previousLoadHead; // @[StoreQueue.scala 103:75:@924.10]
  assign _T_2350 = _T_2348 & _T_2349; // @[StoreQueue.scala 103:49:@925.10]
  assign _T_2352 = _T_2350 == 1'h0; // @[StoreQueue.scala 103:9:@926.10]
  assign _T_2353 = _T_2107 & _T_2352; // @[StoreQueue.scala 102:49:@927.10]
  assign _GEN_720 = _T_2353 ? 1'h0 : checkBits_8; // @[StoreQueue.scala 103:96:@928.10]
  assign _GEN_721 = _T_2345 ? 1'h0 : _GEN_720; // @[StoreQueue.scala 100:102:@918.8]
  assign _GEN_722 = io_loadEmpty ? 1'h0 : _GEN_721; // @[StoreQueue.scala 98:26:@911.6]
  assign _GEN_723 = initBits_8 ? _T_2341 : _GEN_722; // @[StoreQueue.scala 94:35:@896.4]
  assign _T_2366 = _GEN_321 + 4'h1; // @[util.scala 10:8:@939.6]
  assign _GEN_57 = _T_2366 % 5'h10; // @[util.scala 10:14:@940.6]
  assign _T_2367 = _GEN_57[4:0]; // @[util.scala 10:14:@940.6]
  assign _T_2368 = _T_2367 == _GEN_1203; // @[StoreQueue.scala 96:56:@941.6]
  assign _T_2369 = io_loadEmpty & _T_2368; // @[StoreQueue.scala 95:50:@942.6]
  assign _T_2371 = _T_2369 == 1'h0; // @[StoreQueue.scala 95:35:@943.6]
  assign _T_2373 = previousLoadHead <= offsetQ_9; // @[StoreQueue.scala 100:35:@951.8]
  assign _T_2374 = offsetQ_9 < io_loadHead; // @[StoreQueue.scala 100:87:@952.8]
  assign _T_2375 = _T_2373 & _T_2374; // @[StoreQueue.scala 100:61:@953.8]
  assign _T_2378 = io_loadHead <= offsetQ_9; // @[StoreQueue.scala 103:23:@959.10]
  assign _T_2379 = offsetQ_9 < previousLoadHead; // @[StoreQueue.scala 103:75:@960.10]
  assign _T_2380 = _T_2378 & _T_2379; // @[StoreQueue.scala 103:49:@961.10]
  assign _T_2382 = _T_2380 == 1'h0; // @[StoreQueue.scala 103:9:@962.10]
  assign _T_2383 = _T_2107 & _T_2382; // @[StoreQueue.scala 102:49:@963.10]
  assign _GEN_740 = _T_2383 ? 1'h0 : checkBits_9; // @[StoreQueue.scala 103:96:@964.10]
  assign _GEN_741 = _T_2375 ? 1'h0 : _GEN_740; // @[StoreQueue.scala 100:102:@954.8]
  assign _GEN_742 = io_loadEmpty ? 1'h0 : _GEN_741; // @[StoreQueue.scala 98:26:@947.6]
  assign _GEN_743 = initBits_9 ? _T_2371 : _GEN_742; // @[StoreQueue.scala 94:35:@932.4]
  assign _T_2396 = _GEN_355 + 4'h1; // @[util.scala 10:8:@975.6]
  assign _GEN_58 = _T_2396 % 5'h10; // @[util.scala 10:14:@976.6]
  assign _T_2397 = _GEN_58[4:0]; // @[util.scala 10:14:@976.6]
  assign _T_2398 = _T_2397 == _GEN_1203; // @[StoreQueue.scala 96:56:@977.6]
  assign _T_2399 = io_loadEmpty & _T_2398; // @[StoreQueue.scala 95:50:@978.6]
  assign _T_2401 = _T_2399 == 1'h0; // @[StoreQueue.scala 95:35:@979.6]
  assign _T_2403 = previousLoadHead <= offsetQ_10; // @[StoreQueue.scala 100:35:@987.8]
  assign _T_2404 = offsetQ_10 < io_loadHead; // @[StoreQueue.scala 100:87:@988.8]
  assign _T_2405 = _T_2403 & _T_2404; // @[StoreQueue.scala 100:61:@989.8]
  assign _T_2408 = io_loadHead <= offsetQ_10; // @[StoreQueue.scala 103:23:@995.10]
  assign _T_2409 = offsetQ_10 < previousLoadHead; // @[StoreQueue.scala 103:75:@996.10]
  assign _T_2410 = _T_2408 & _T_2409; // @[StoreQueue.scala 103:49:@997.10]
  assign _T_2412 = _T_2410 == 1'h0; // @[StoreQueue.scala 103:9:@998.10]
  assign _T_2413 = _T_2107 & _T_2412; // @[StoreQueue.scala 102:49:@999.10]
  assign _GEN_760 = _T_2413 ? 1'h0 : checkBits_10; // @[StoreQueue.scala 103:96:@1000.10]
  assign _GEN_761 = _T_2405 ? 1'h0 : _GEN_760; // @[StoreQueue.scala 100:102:@990.8]
  assign _GEN_762 = io_loadEmpty ? 1'h0 : _GEN_761; // @[StoreQueue.scala 98:26:@983.6]
  assign _GEN_763 = initBits_10 ? _T_2401 : _GEN_762; // @[StoreQueue.scala 94:35:@968.4]
  assign _T_2426 = _GEN_389 + 4'h1; // @[util.scala 10:8:@1011.6]
  assign _GEN_59 = _T_2426 % 5'h10; // @[util.scala 10:14:@1012.6]
  assign _T_2427 = _GEN_59[4:0]; // @[util.scala 10:14:@1012.6]
  assign _T_2428 = _T_2427 == _GEN_1203; // @[StoreQueue.scala 96:56:@1013.6]
  assign _T_2429 = io_loadEmpty & _T_2428; // @[StoreQueue.scala 95:50:@1014.6]
  assign _T_2431 = _T_2429 == 1'h0; // @[StoreQueue.scala 95:35:@1015.6]
  assign _T_2433 = previousLoadHead <= offsetQ_11; // @[StoreQueue.scala 100:35:@1023.8]
  assign _T_2434 = offsetQ_11 < io_loadHead; // @[StoreQueue.scala 100:87:@1024.8]
  assign _T_2435 = _T_2433 & _T_2434; // @[StoreQueue.scala 100:61:@1025.8]
  assign _T_2438 = io_loadHead <= offsetQ_11; // @[StoreQueue.scala 103:23:@1031.10]
  assign _T_2439 = offsetQ_11 < previousLoadHead; // @[StoreQueue.scala 103:75:@1032.10]
  assign _T_2440 = _T_2438 & _T_2439; // @[StoreQueue.scala 103:49:@1033.10]
  assign _T_2442 = _T_2440 == 1'h0; // @[StoreQueue.scala 103:9:@1034.10]
  assign _T_2443 = _T_2107 & _T_2442; // @[StoreQueue.scala 102:49:@1035.10]
  assign _GEN_780 = _T_2443 ? 1'h0 : checkBits_11; // @[StoreQueue.scala 103:96:@1036.10]
  assign _GEN_781 = _T_2435 ? 1'h0 : _GEN_780; // @[StoreQueue.scala 100:102:@1026.8]
  assign _GEN_782 = io_loadEmpty ? 1'h0 : _GEN_781; // @[StoreQueue.scala 98:26:@1019.6]
  assign _GEN_783 = initBits_11 ? _T_2431 : _GEN_782; // @[StoreQueue.scala 94:35:@1004.4]
  assign _T_2456 = _GEN_423 + 4'h1; // @[util.scala 10:8:@1047.6]
  assign _GEN_60 = _T_2456 % 5'h10; // @[util.scala 10:14:@1048.6]
  assign _T_2457 = _GEN_60[4:0]; // @[util.scala 10:14:@1048.6]
  assign _T_2458 = _T_2457 == _GEN_1203; // @[StoreQueue.scala 96:56:@1049.6]
  assign _T_2459 = io_loadEmpty & _T_2458; // @[StoreQueue.scala 95:50:@1050.6]
  assign _T_2461 = _T_2459 == 1'h0; // @[StoreQueue.scala 95:35:@1051.6]
  assign _T_2463 = previousLoadHead <= offsetQ_12; // @[StoreQueue.scala 100:35:@1059.8]
  assign _T_2464 = offsetQ_12 < io_loadHead; // @[StoreQueue.scala 100:87:@1060.8]
  assign _T_2465 = _T_2463 & _T_2464; // @[StoreQueue.scala 100:61:@1061.8]
  assign _T_2468 = io_loadHead <= offsetQ_12; // @[StoreQueue.scala 103:23:@1067.10]
  assign _T_2469 = offsetQ_12 < previousLoadHead; // @[StoreQueue.scala 103:75:@1068.10]
  assign _T_2470 = _T_2468 & _T_2469; // @[StoreQueue.scala 103:49:@1069.10]
  assign _T_2472 = _T_2470 == 1'h0; // @[StoreQueue.scala 103:9:@1070.10]
  assign _T_2473 = _T_2107 & _T_2472; // @[StoreQueue.scala 102:49:@1071.10]
  assign _GEN_800 = _T_2473 ? 1'h0 : checkBits_12; // @[StoreQueue.scala 103:96:@1072.10]
  assign _GEN_801 = _T_2465 ? 1'h0 : _GEN_800; // @[StoreQueue.scala 100:102:@1062.8]
  assign _GEN_802 = io_loadEmpty ? 1'h0 : _GEN_801; // @[StoreQueue.scala 98:26:@1055.6]
  assign _GEN_803 = initBits_12 ? _T_2461 : _GEN_802; // @[StoreQueue.scala 94:35:@1040.4]
  assign _T_2486 = _GEN_457 + 4'h1; // @[util.scala 10:8:@1083.6]
  assign _GEN_61 = _T_2486 % 5'h10; // @[util.scala 10:14:@1084.6]
  assign _T_2487 = _GEN_61[4:0]; // @[util.scala 10:14:@1084.6]
  assign _T_2488 = _T_2487 == _GEN_1203; // @[StoreQueue.scala 96:56:@1085.6]
  assign _T_2489 = io_loadEmpty & _T_2488; // @[StoreQueue.scala 95:50:@1086.6]
  assign _T_2491 = _T_2489 == 1'h0; // @[StoreQueue.scala 95:35:@1087.6]
  assign _T_2493 = previousLoadHead <= offsetQ_13; // @[StoreQueue.scala 100:35:@1095.8]
  assign _T_2494 = offsetQ_13 < io_loadHead; // @[StoreQueue.scala 100:87:@1096.8]
  assign _T_2495 = _T_2493 & _T_2494; // @[StoreQueue.scala 100:61:@1097.8]
  assign _T_2498 = io_loadHead <= offsetQ_13; // @[StoreQueue.scala 103:23:@1103.10]
  assign _T_2499 = offsetQ_13 < previousLoadHead; // @[StoreQueue.scala 103:75:@1104.10]
  assign _T_2500 = _T_2498 & _T_2499; // @[StoreQueue.scala 103:49:@1105.10]
  assign _T_2502 = _T_2500 == 1'h0; // @[StoreQueue.scala 103:9:@1106.10]
  assign _T_2503 = _T_2107 & _T_2502; // @[StoreQueue.scala 102:49:@1107.10]
  assign _GEN_820 = _T_2503 ? 1'h0 : checkBits_13; // @[StoreQueue.scala 103:96:@1108.10]
  assign _GEN_821 = _T_2495 ? 1'h0 : _GEN_820; // @[StoreQueue.scala 100:102:@1098.8]
  assign _GEN_822 = io_loadEmpty ? 1'h0 : _GEN_821; // @[StoreQueue.scala 98:26:@1091.6]
  assign _GEN_823 = initBits_13 ? _T_2491 : _GEN_822; // @[StoreQueue.scala 94:35:@1076.4]
  assign _T_2516 = _GEN_491 + 4'h1; // @[util.scala 10:8:@1119.6]
  assign _GEN_62 = _T_2516 % 5'h10; // @[util.scala 10:14:@1120.6]
  assign _T_2517 = _GEN_62[4:0]; // @[util.scala 10:14:@1120.6]
  assign _T_2518 = _T_2517 == _GEN_1203; // @[StoreQueue.scala 96:56:@1121.6]
  assign _T_2519 = io_loadEmpty & _T_2518; // @[StoreQueue.scala 95:50:@1122.6]
  assign _T_2521 = _T_2519 == 1'h0; // @[StoreQueue.scala 95:35:@1123.6]
  assign _T_2523 = previousLoadHead <= offsetQ_14; // @[StoreQueue.scala 100:35:@1131.8]
  assign _T_2524 = offsetQ_14 < io_loadHead; // @[StoreQueue.scala 100:87:@1132.8]
  assign _T_2525 = _T_2523 & _T_2524; // @[StoreQueue.scala 100:61:@1133.8]
  assign _T_2528 = io_loadHead <= offsetQ_14; // @[StoreQueue.scala 103:23:@1139.10]
  assign _T_2529 = offsetQ_14 < previousLoadHead; // @[StoreQueue.scala 103:75:@1140.10]
  assign _T_2530 = _T_2528 & _T_2529; // @[StoreQueue.scala 103:49:@1141.10]
  assign _T_2532 = _T_2530 == 1'h0; // @[StoreQueue.scala 103:9:@1142.10]
  assign _T_2533 = _T_2107 & _T_2532; // @[StoreQueue.scala 102:49:@1143.10]
  assign _GEN_840 = _T_2533 ? 1'h0 : checkBits_14; // @[StoreQueue.scala 103:96:@1144.10]
  assign _GEN_841 = _T_2525 ? 1'h0 : _GEN_840; // @[StoreQueue.scala 100:102:@1134.8]
  assign _GEN_842 = io_loadEmpty ? 1'h0 : _GEN_841; // @[StoreQueue.scala 98:26:@1127.6]
  assign _GEN_843 = initBits_14 ? _T_2521 : _GEN_842; // @[StoreQueue.scala 94:35:@1112.4]
  assign _T_2546 = _GEN_525 + 4'h1; // @[util.scala 10:8:@1155.6]
  assign _GEN_63 = _T_2546 % 5'h10; // @[util.scala 10:14:@1156.6]
  assign _T_2547 = _GEN_63[4:0]; // @[util.scala 10:14:@1156.6]
  assign _T_2548 = _T_2547 == _GEN_1203; // @[StoreQueue.scala 96:56:@1157.6]
  assign _T_2549 = io_loadEmpty & _T_2548; // @[StoreQueue.scala 95:50:@1158.6]
  assign _T_2551 = _T_2549 == 1'h0; // @[StoreQueue.scala 95:35:@1159.6]
  assign _T_2553 = previousLoadHead <= offsetQ_15; // @[StoreQueue.scala 100:35:@1167.8]
  assign _T_2554 = offsetQ_15 < io_loadHead; // @[StoreQueue.scala 100:87:@1168.8]
  assign _T_2555 = _T_2553 & _T_2554; // @[StoreQueue.scala 100:61:@1169.8]
  assign _T_2558 = io_loadHead <= offsetQ_15; // @[StoreQueue.scala 103:23:@1175.10]
  assign _T_2559 = offsetQ_15 < previousLoadHead; // @[StoreQueue.scala 103:75:@1176.10]
  assign _T_2560 = _T_2558 & _T_2559; // @[StoreQueue.scala 103:49:@1177.10]
  assign _T_2562 = _T_2560 == 1'h0; // @[StoreQueue.scala 103:9:@1178.10]
  assign _T_2563 = _T_2107 & _T_2562; // @[StoreQueue.scala 102:49:@1179.10]
  assign _GEN_860 = _T_2563 ? 1'h0 : checkBits_15; // @[StoreQueue.scala 103:96:@1180.10]
  assign _GEN_861 = _T_2555 ? 1'h0 : _GEN_860; // @[StoreQueue.scala 100:102:@1170.8]
  assign _GEN_862 = io_loadEmpty ? 1'h0 : _GEN_861; // @[StoreQueue.scala 98:26:@1163.6]
  assign _GEN_863 = initBits_15 ? _T_2551 : _GEN_862; // @[StoreQueue.scala 94:35:@1148.4]
  assign _T_2565 = io_loadHead < io_loadTail; // @[StoreQueue.scala 119:103:@1184.4]
  assign _T_2567 = io_loadHead <= 4'h0; // @[StoreQueue.scala 120:17:@1185.4]
  assign _T_2569 = 4'h0 < io_loadTail; // @[StoreQueue.scala 120:35:@1186.4]
  assign _T_2570 = _T_2567 & _T_2569; // @[StoreQueue.scala 120:26:@1187.4]
  assign _T_2572 = io_loadEmpty == 1'h0; // @[StoreQueue.scala 120:50:@1188.4]
  assign _T_2574 = io_loadTail <= 4'h0; // @[StoreQueue.scala 120:81:@1189.4]
  assign _T_2576 = 4'h0 < io_loadHead; // @[StoreQueue.scala 120:99:@1190.4]
  assign _T_2577 = _T_2574 & _T_2576; // @[StoreQueue.scala 120:90:@1191.4]
  assign _T_2579 = _T_2577 == 1'h0; // @[StoreQueue.scala 120:67:@1192.4]
  assign _T_2580 = _T_2572 & _T_2579; // @[StoreQueue.scala 120:64:@1193.4]
  assign validEntriesInLoadQ_0 = _T_2565 ? _T_2570 : _T_2580; // @[StoreQueue.scala 119:90:@1194.4]
  assign _T_2584 = io_loadHead <= 4'h1; // @[StoreQueue.scala 120:17:@1196.4]
  assign _T_2586 = 4'h1 < io_loadTail; // @[StoreQueue.scala 120:35:@1197.4]
  assign _T_2587 = _T_2584 & _T_2586; // @[StoreQueue.scala 120:26:@1198.4]
  assign _T_2591 = io_loadTail <= 4'h1; // @[StoreQueue.scala 120:81:@1200.4]
  assign _T_2593 = 4'h1 < io_loadHead; // @[StoreQueue.scala 120:99:@1201.4]
  assign _T_2594 = _T_2591 & _T_2593; // @[StoreQueue.scala 120:90:@1202.4]
  assign _T_2596 = _T_2594 == 1'h0; // @[StoreQueue.scala 120:67:@1203.4]
  assign _T_2597 = _T_2572 & _T_2596; // @[StoreQueue.scala 120:64:@1204.4]
  assign validEntriesInLoadQ_1 = _T_2565 ? _T_2587 : _T_2597; // @[StoreQueue.scala 119:90:@1205.4]
  assign _T_2601 = io_loadHead <= 4'h2; // @[StoreQueue.scala 120:17:@1207.4]
  assign _T_2603 = 4'h2 < io_loadTail; // @[StoreQueue.scala 120:35:@1208.4]
  assign _T_2604 = _T_2601 & _T_2603; // @[StoreQueue.scala 120:26:@1209.4]
  assign _T_2608 = io_loadTail <= 4'h2; // @[StoreQueue.scala 120:81:@1211.4]
  assign _T_2610 = 4'h2 < io_loadHead; // @[StoreQueue.scala 120:99:@1212.4]
  assign _T_2611 = _T_2608 & _T_2610; // @[StoreQueue.scala 120:90:@1213.4]
  assign _T_2613 = _T_2611 == 1'h0; // @[StoreQueue.scala 120:67:@1214.4]
  assign _T_2614 = _T_2572 & _T_2613; // @[StoreQueue.scala 120:64:@1215.4]
  assign validEntriesInLoadQ_2 = _T_2565 ? _T_2604 : _T_2614; // @[StoreQueue.scala 119:90:@1216.4]
  assign _T_2618 = io_loadHead <= 4'h3; // @[StoreQueue.scala 120:17:@1218.4]
  assign _T_2620 = 4'h3 < io_loadTail; // @[StoreQueue.scala 120:35:@1219.4]
  assign _T_2621 = _T_2618 & _T_2620; // @[StoreQueue.scala 120:26:@1220.4]
  assign _T_2625 = io_loadTail <= 4'h3; // @[StoreQueue.scala 120:81:@1222.4]
  assign _T_2627 = 4'h3 < io_loadHead; // @[StoreQueue.scala 120:99:@1223.4]
  assign _T_2628 = _T_2625 & _T_2627; // @[StoreQueue.scala 120:90:@1224.4]
  assign _T_2630 = _T_2628 == 1'h0; // @[StoreQueue.scala 120:67:@1225.4]
  assign _T_2631 = _T_2572 & _T_2630; // @[StoreQueue.scala 120:64:@1226.4]
  assign validEntriesInLoadQ_3 = _T_2565 ? _T_2621 : _T_2631; // @[StoreQueue.scala 119:90:@1227.4]
  assign _T_2635 = io_loadHead <= 4'h4; // @[StoreQueue.scala 120:17:@1229.4]
  assign _T_2637 = 4'h4 < io_loadTail; // @[StoreQueue.scala 120:35:@1230.4]
  assign _T_2638 = _T_2635 & _T_2637; // @[StoreQueue.scala 120:26:@1231.4]
  assign _T_2642 = io_loadTail <= 4'h4; // @[StoreQueue.scala 120:81:@1233.4]
  assign _T_2644 = 4'h4 < io_loadHead; // @[StoreQueue.scala 120:99:@1234.4]
  assign _T_2645 = _T_2642 & _T_2644; // @[StoreQueue.scala 120:90:@1235.4]
  assign _T_2647 = _T_2645 == 1'h0; // @[StoreQueue.scala 120:67:@1236.4]
  assign _T_2648 = _T_2572 & _T_2647; // @[StoreQueue.scala 120:64:@1237.4]
  assign validEntriesInLoadQ_4 = _T_2565 ? _T_2638 : _T_2648; // @[StoreQueue.scala 119:90:@1238.4]
  assign _T_2652 = io_loadHead <= 4'h5; // @[StoreQueue.scala 120:17:@1240.4]
  assign _T_2654 = 4'h5 < io_loadTail; // @[StoreQueue.scala 120:35:@1241.4]
  assign _T_2655 = _T_2652 & _T_2654; // @[StoreQueue.scala 120:26:@1242.4]
  assign _T_2659 = io_loadTail <= 4'h5; // @[StoreQueue.scala 120:81:@1244.4]
  assign _T_2661 = 4'h5 < io_loadHead; // @[StoreQueue.scala 120:99:@1245.4]
  assign _T_2662 = _T_2659 & _T_2661; // @[StoreQueue.scala 120:90:@1246.4]
  assign _T_2664 = _T_2662 == 1'h0; // @[StoreQueue.scala 120:67:@1247.4]
  assign _T_2665 = _T_2572 & _T_2664; // @[StoreQueue.scala 120:64:@1248.4]
  assign validEntriesInLoadQ_5 = _T_2565 ? _T_2655 : _T_2665; // @[StoreQueue.scala 119:90:@1249.4]
  assign _T_2669 = io_loadHead <= 4'h6; // @[StoreQueue.scala 120:17:@1251.4]
  assign _T_2671 = 4'h6 < io_loadTail; // @[StoreQueue.scala 120:35:@1252.4]
  assign _T_2672 = _T_2669 & _T_2671; // @[StoreQueue.scala 120:26:@1253.4]
  assign _T_2676 = io_loadTail <= 4'h6; // @[StoreQueue.scala 120:81:@1255.4]
  assign _T_2678 = 4'h6 < io_loadHead; // @[StoreQueue.scala 120:99:@1256.4]
  assign _T_2679 = _T_2676 & _T_2678; // @[StoreQueue.scala 120:90:@1257.4]
  assign _T_2681 = _T_2679 == 1'h0; // @[StoreQueue.scala 120:67:@1258.4]
  assign _T_2682 = _T_2572 & _T_2681; // @[StoreQueue.scala 120:64:@1259.4]
  assign validEntriesInLoadQ_6 = _T_2565 ? _T_2672 : _T_2682; // @[StoreQueue.scala 119:90:@1260.4]
  assign _T_2686 = io_loadHead <= 4'h7; // @[StoreQueue.scala 120:17:@1262.4]
  assign _T_2688 = 4'h7 < io_loadTail; // @[StoreQueue.scala 120:35:@1263.4]
  assign _T_2689 = _T_2686 & _T_2688; // @[StoreQueue.scala 120:26:@1264.4]
  assign _T_2693 = io_loadTail <= 4'h7; // @[StoreQueue.scala 120:81:@1266.4]
  assign _T_2695 = 4'h7 < io_loadHead; // @[StoreQueue.scala 120:99:@1267.4]
  assign _T_2696 = _T_2693 & _T_2695; // @[StoreQueue.scala 120:90:@1268.4]
  assign _T_2698 = _T_2696 == 1'h0; // @[StoreQueue.scala 120:67:@1269.4]
  assign _T_2699 = _T_2572 & _T_2698; // @[StoreQueue.scala 120:64:@1270.4]
  assign validEntriesInLoadQ_7 = _T_2565 ? _T_2689 : _T_2699; // @[StoreQueue.scala 119:90:@1271.4]
  assign _T_2703 = io_loadHead <= 4'h8; // @[StoreQueue.scala 120:17:@1273.4]
  assign _T_2705 = 4'h8 < io_loadTail; // @[StoreQueue.scala 120:35:@1274.4]
  assign _T_2706 = _T_2703 & _T_2705; // @[StoreQueue.scala 120:26:@1275.4]
  assign _T_2710 = io_loadTail <= 4'h8; // @[StoreQueue.scala 120:81:@1277.4]
  assign _T_2712 = 4'h8 < io_loadHead; // @[StoreQueue.scala 120:99:@1278.4]
  assign _T_2713 = _T_2710 & _T_2712; // @[StoreQueue.scala 120:90:@1279.4]
  assign _T_2715 = _T_2713 == 1'h0; // @[StoreQueue.scala 120:67:@1280.4]
  assign _T_2716 = _T_2572 & _T_2715; // @[StoreQueue.scala 120:64:@1281.4]
  assign validEntriesInLoadQ_8 = _T_2565 ? _T_2706 : _T_2716; // @[StoreQueue.scala 119:90:@1282.4]
  assign _T_2720 = io_loadHead <= 4'h9; // @[StoreQueue.scala 120:17:@1284.4]
  assign _T_2722 = 4'h9 < io_loadTail; // @[StoreQueue.scala 120:35:@1285.4]
  assign _T_2723 = _T_2720 & _T_2722; // @[StoreQueue.scala 120:26:@1286.4]
  assign _T_2727 = io_loadTail <= 4'h9; // @[StoreQueue.scala 120:81:@1288.4]
  assign _T_2729 = 4'h9 < io_loadHead; // @[StoreQueue.scala 120:99:@1289.4]
  assign _T_2730 = _T_2727 & _T_2729; // @[StoreQueue.scala 120:90:@1290.4]
  assign _T_2732 = _T_2730 == 1'h0; // @[StoreQueue.scala 120:67:@1291.4]
  assign _T_2733 = _T_2572 & _T_2732; // @[StoreQueue.scala 120:64:@1292.4]
  assign validEntriesInLoadQ_9 = _T_2565 ? _T_2723 : _T_2733; // @[StoreQueue.scala 119:90:@1293.4]
  assign _T_2737 = io_loadHead <= 4'ha; // @[StoreQueue.scala 120:17:@1295.4]
  assign _T_2739 = 4'ha < io_loadTail; // @[StoreQueue.scala 120:35:@1296.4]
  assign _T_2740 = _T_2737 & _T_2739; // @[StoreQueue.scala 120:26:@1297.4]
  assign _T_2744 = io_loadTail <= 4'ha; // @[StoreQueue.scala 120:81:@1299.4]
  assign _T_2746 = 4'ha < io_loadHead; // @[StoreQueue.scala 120:99:@1300.4]
  assign _T_2747 = _T_2744 & _T_2746; // @[StoreQueue.scala 120:90:@1301.4]
  assign _T_2749 = _T_2747 == 1'h0; // @[StoreQueue.scala 120:67:@1302.4]
  assign _T_2750 = _T_2572 & _T_2749; // @[StoreQueue.scala 120:64:@1303.4]
  assign validEntriesInLoadQ_10 = _T_2565 ? _T_2740 : _T_2750; // @[StoreQueue.scala 119:90:@1304.4]
  assign _T_2754 = io_loadHead <= 4'hb; // @[StoreQueue.scala 120:17:@1306.4]
  assign _T_2756 = 4'hb < io_loadTail; // @[StoreQueue.scala 120:35:@1307.4]
  assign _T_2757 = _T_2754 & _T_2756; // @[StoreQueue.scala 120:26:@1308.4]
  assign _T_2761 = io_loadTail <= 4'hb; // @[StoreQueue.scala 120:81:@1310.4]
  assign _T_2763 = 4'hb < io_loadHead; // @[StoreQueue.scala 120:99:@1311.4]
  assign _T_2764 = _T_2761 & _T_2763; // @[StoreQueue.scala 120:90:@1312.4]
  assign _T_2766 = _T_2764 == 1'h0; // @[StoreQueue.scala 120:67:@1313.4]
  assign _T_2767 = _T_2572 & _T_2766; // @[StoreQueue.scala 120:64:@1314.4]
  assign validEntriesInLoadQ_11 = _T_2565 ? _T_2757 : _T_2767; // @[StoreQueue.scala 119:90:@1315.4]
  assign _T_2771 = io_loadHead <= 4'hc; // @[StoreQueue.scala 120:17:@1317.4]
  assign _T_2773 = 4'hc < io_loadTail; // @[StoreQueue.scala 120:35:@1318.4]
  assign _T_2774 = _T_2771 & _T_2773; // @[StoreQueue.scala 120:26:@1319.4]
  assign _T_2778 = io_loadTail <= 4'hc; // @[StoreQueue.scala 120:81:@1321.4]
  assign _T_2780 = 4'hc < io_loadHead; // @[StoreQueue.scala 120:99:@1322.4]
  assign _T_2781 = _T_2778 & _T_2780; // @[StoreQueue.scala 120:90:@1323.4]
  assign _T_2783 = _T_2781 == 1'h0; // @[StoreQueue.scala 120:67:@1324.4]
  assign _T_2784 = _T_2572 & _T_2783; // @[StoreQueue.scala 120:64:@1325.4]
  assign validEntriesInLoadQ_12 = _T_2565 ? _T_2774 : _T_2784; // @[StoreQueue.scala 119:90:@1326.4]
  assign _T_2788 = io_loadHead <= 4'hd; // @[StoreQueue.scala 120:17:@1328.4]
  assign _T_2790 = 4'hd < io_loadTail; // @[StoreQueue.scala 120:35:@1329.4]
  assign _T_2791 = _T_2788 & _T_2790; // @[StoreQueue.scala 120:26:@1330.4]
  assign _T_2795 = io_loadTail <= 4'hd; // @[StoreQueue.scala 120:81:@1332.4]
  assign _T_2797 = 4'hd < io_loadHead; // @[StoreQueue.scala 120:99:@1333.4]
  assign _T_2798 = _T_2795 & _T_2797; // @[StoreQueue.scala 120:90:@1334.4]
  assign _T_2800 = _T_2798 == 1'h0; // @[StoreQueue.scala 120:67:@1335.4]
  assign _T_2801 = _T_2572 & _T_2800; // @[StoreQueue.scala 120:64:@1336.4]
  assign validEntriesInLoadQ_13 = _T_2565 ? _T_2791 : _T_2801; // @[StoreQueue.scala 119:90:@1337.4]
  assign _T_2805 = io_loadHead <= 4'he; // @[StoreQueue.scala 120:17:@1339.4]
  assign _T_2807 = 4'he < io_loadTail; // @[StoreQueue.scala 120:35:@1340.4]
  assign _T_2808 = _T_2805 & _T_2807; // @[StoreQueue.scala 120:26:@1341.4]
  assign _T_2812 = io_loadTail <= 4'he; // @[StoreQueue.scala 120:81:@1343.4]
  assign _T_2814 = 4'he < io_loadHead; // @[StoreQueue.scala 120:99:@1344.4]
  assign _T_2815 = _T_2812 & _T_2814; // @[StoreQueue.scala 120:90:@1345.4]
  assign _T_2817 = _T_2815 == 1'h0; // @[StoreQueue.scala 120:67:@1346.4]
  assign _T_2818 = _T_2572 & _T_2817; // @[StoreQueue.scala 120:64:@1347.4]
  assign validEntriesInLoadQ_14 = _T_2565 ? _T_2808 : _T_2818; // @[StoreQueue.scala 119:90:@1348.4]
  assign validEntriesInLoadQ_15 = _T_2565 ? 1'h0 : _T_2572; // @[StoreQueue.scala 119:90:@1359.4]
  assign _GEN_865 = 4'h1 == head ? offsetQ_1 : offsetQ_0; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_866 = 4'h2 == head ? offsetQ_2 : _GEN_865; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_867 = 4'h3 == head ? offsetQ_3 : _GEN_866; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_868 = 4'h4 == head ? offsetQ_4 : _GEN_867; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_869 = 4'h5 == head ? offsetQ_5 : _GEN_868; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_870 = 4'h6 == head ? offsetQ_6 : _GEN_869; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_871 = 4'h7 == head ? offsetQ_7 : _GEN_870; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_872 = 4'h8 == head ? offsetQ_8 : _GEN_871; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_873 = 4'h9 == head ? offsetQ_9 : _GEN_872; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_874 = 4'ha == head ? offsetQ_10 : _GEN_873; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_875 = 4'hb == head ? offsetQ_11 : _GEN_874; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_876 = 4'hc == head ? offsetQ_12 : _GEN_875; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_877 = 4'hd == head ? offsetQ_13 : _GEN_876; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_878 = 4'he == head ? offsetQ_14 : _GEN_877; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_879 = 4'hf == head ? offsetQ_15 : _GEN_878; // @[StoreQueue.scala 126:96:@1377.4]
  assign _T_2861 = io_loadHead <= _GEN_879; // @[StoreQueue.scala 126:96:@1377.4]
  assign loadsToCheck_0 = _T_2861 ? _T_2567 : 1'h1; // @[StoreQueue.scala 126:83:@1385.4]
  assign _T_2891 = 4'h1 <= _GEN_879; // @[StoreQueue.scala 127:37:@1388.4]
  assign _T_2892 = _T_2584 & _T_2891; // @[StoreQueue.scala 127:28:@1389.4]
  assign _T_2897 = _GEN_879 < 4'h1; // @[StoreQueue.scala 127:71:@1390.4]
  assign _T_2900 = _T_2897 & _T_2593; // @[StoreQueue.scala 127:79:@1392.4]
  assign _T_2902 = _T_2900 == 1'h0; // @[StoreQueue.scala 127:55:@1393.4]
  assign loadsToCheck_1 = _T_2861 ? _T_2892 : _T_2902; // @[StoreQueue.scala 126:83:@1394.4]
  assign _T_2914 = 4'h2 <= _GEN_879; // @[StoreQueue.scala 127:37:@1397.4]
  assign _T_2915 = _T_2601 & _T_2914; // @[StoreQueue.scala 127:28:@1398.4]
  assign _T_2920 = _GEN_879 < 4'h2; // @[StoreQueue.scala 127:71:@1399.4]
  assign _T_2923 = _T_2920 & _T_2610; // @[StoreQueue.scala 127:79:@1401.4]
  assign _T_2925 = _T_2923 == 1'h0; // @[StoreQueue.scala 127:55:@1402.4]
  assign loadsToCheck_2 = _T_2861 ? _T_2915 : _T_2925; // @[StoreQueue.scala 126:83:@1403.4]
  assign _T_2937 = 4'h3 <= _GEN_879; // @[StoreQueue.scala 127:37:@1406.4]
  assign _T_2938 = _T_2618 & _T_2937; // @[StoreQueue.scala 127:28:@1407.4]
  assign _T_2943 = _GEN_879 < 4'h3; // @[StoreQueue.scala 127:71:@1408.4]
  assign _T_2946 = _T_2943 & _T_2627; // @[StoreQueue.scala 127:79:@1410.4]
  assign _T_2948 = _T_2946 == 1'h0; // @[StoreQueue.scala 127:55:@1411.4]
  assign loadsToCheck_3 = _T_2861 ? _T_2938 : _T_2948; // @[StoreQueue.scala 126:83:@1412.4]
  assign _T_2960 = 4'h4 <= _GEN_879; // @[StoreQueue.scala 127:37:@1415.4]
  assign _T_2961 = _T_2635 & _T_2960; // @[StoreQueue.scala 127:28:@1416.4]
  assign _T_2966 = _GEN_879 < 4'h4; // @[StoreQueue.scala 127:71:@1417.4]
  assign _T_2969 = _T_2966 & _T_2644; // @[StoreQueue.scala 127:79:@1419.4]
  assign _T_2971 = _T_2969 == 1'h0; // @[StoreQueue.scala 127:55:@1420.4]
  assign loadsToCheck_4 = _T_2861 ? _T_2961 : _T_2971; // @[StoreQueue.scala 126:83:@1421.4]
  assign _T_2983 = 4'h5 <= _GEN_879; // @[StoreQueue.scala 127:37:@1424.4]
  assign _T_2984 = _T_2652 & _T_2983; // @[StoreQueue.scala 127:28:@1425.4]
  assign _T_2989 = _GEN_879 < 4'h5; // @[StoreQueue.scala 127:71:@1426.4]
  assign _T_2992 = _T_2989 & _T_2661; // @[StoreQueue.scala 127:79:@1428.4]
  assign _T_2994 = _T_2992 == 1'h0; // @[StoreQueue.scala 127:55:@1429.4]
  assign loadsToCheck_5 = _T_2861 ? _T_2984 : _T_2994; // @[StoreQueue.scala 126:83:@1430.4]
  assign _T_3006 = 4'h6 <= _GEN_879; // @[StoreQueue.scala 127:37:@1433.4]
  assign _T_3007 = _T_2669 & _T_3006; // @[StoreQueue.scala 127:28:@1434.4]
  assign _T_3012 = _GEN_879 < 4'h6; // @[StoreQueue.scala 127:71:@1435.4]
  assign _T_3015 = _T_3012 & _T_2678; // @[StoreQueue.scala 127:79:@1437.4]
  assign _T_3017 = _T_3015 == 1'h0; // @[StoreQueue.scala 127:55:@1438.4]
  assign loadsToCheck_6 = _T_2861 ? _T_3007 : _T_3017; // @[StoreQueue.scala 126:83:@1439.4]
  assign _T_3029 = 4'h7 <= _GEN_879; // @[StoreQueue.scala 127:37:@1442.4]
  assign _T_3030 = _T_2686 & _T_3029; // @[StoreQueue.scala 127:28:@1443.4]
  assign _T_3035 = _GEN_879 < 4'h7; // @[StoreQueue.scala 127:71:@1444.4]
  assign _T_3038 = _T_3035 & _T_2695; // @[StoreQueue.scala 127:79:@1446.4]
  assign _T_3040 = _T_3038 == 1'h0; // @[StoreQueue.scala 127:55:@1447.4]
  assign loadsToCheck_7 = _T_2861 ? _T_3030 : _T_3040; // @[StoreQueue.scala 126:83:@1448.4]
  assign _T_3052 = 4'h8 <= _GEN_879; // @[StoreQueue.scala 127:37:@1451.4]
  assign _T_3053 = _T_2703 & _T_3052; // @[StoreQueue.scala 127:28:@1452.4]
  assign _T_3058 = _GEN_879 < 4'h8; // @[StoreQueue.scala 127:71:@1453.4]
  assign _T_3061 = _T_3058 & _T_2712; // @[StoreQueue.scala 127:79:@1455.4]
  assign _T_3063 = _T_3061 == 1'h0; // @[StoreQueue.scala 127:55:@1456.4]
  assign loadsToCheck_8 = _T_2861 ? _T_3053 : _T_3063; // @[StoreQueue.scala 126:83:@1457.4]
  assign _T_3075 = 4'h9 <= _GEN_879; // @[StoreQueue.scala 127:37:@1460.4]
  assign _T_3076 = _T_2720 & _T_3075; // @[StoreQueue.scala 127:28:@1461.4]
  assign _T_3081 = _GEN_879 < 4'h9; // @[StoreQueue.scala 127:71:@1462.4]
  assign _T_3084 = _T_3081 & _T_2729; // @[StoreQueue.scala 127:79:@1464.4]
  assign _T_3086 = _T_3084 == 1'h0; // @[StoreQueue.scala 127:55:@1465.4]
  assign loadsToCheck_9 = _T_2861 ? _T_3076 : _T_3086; // @[StoreQueue.scala 126:83:@1466.4]
  assign _T_3098 = 4'ha <= _GEN_879; // @[StoreQueue.scala 127:37:@1469.4]
  assign _T_3099 = _T_2737 & _T_3098; // @[StoreQueue.scala 127:28:@1470.4]
  assign _T_3104 = _GEN_879 < 4'ha; // @[StoreQueue.scala 127:71:@1471.4]
  assign _T_3107 = _T_3104 & _T_2746; // @[StoreQueue.scala 127:79:@1473.4]
  assign _T_3109 = _T_3107 == 1'h0; // @[StoreQueue.scala 127:55:@1474.4]
  assign loadsToCheck_10 = _T_2861 ? _T_3099 : _T_3109; // @[StoreQueue.scala 126:83:@1475.4]
  assign _T_3121 = 4'hb <= _GEN_879; // @[StoreQueue.scala 127:37:@1478.4]
  assign _T_3122 = _T_2754 & _T_3121; // @[StoreQueue.scala 127:28:@1479.4]
  assign _T_3127 = _GEN_879 < 4'hb; // @[StoreQueue.scala 127:71:@1480.4]
  assign _T_3130 = _T_3127 & _T_2763; // @[StoreQueue.scala 127:79:@1482.4]
  assign _T_3132 = _T_3130 == 1'h0; // @[StoreQueue.scala 127:55:@1483.4]
  assign loadsToCheck_11 = _T_2861 ? _T_3122 : _T_3132; // @[StoreQueue.scala 126:83:@1484.4]
  assign _T_3144 = 4'hc <= _GEN_879; // @[StoreQueue.scala 127:37:@1487.4]
  assign _T_3145 = _T_2771 & _T_3144; // @[StoreQueue.scala 127:28:@1488.4]
  assign _T_3150 = _GEN_879 < 4'hc; // @[StoreQueue.scala 127:71:@1489.4]
  assign _T_3153 = _T_3150 & _T_2780; // @[StoreQueue.scala 127:79:@1491.4]
  assign _T_3155 = _T_3153 == 1'h0; // @[StoreQueue.scala 127:55:@1492.4]
  assign loadsToCheck_12 = _T_2861 ? _T_3145 : _T_3155; // @[StoreQueue.scala 126:83:@1493.4]
  assign _T_3167 = 4'hd <= _GEN_879; // @[StoreQueue.scala 127:37:@1496.4]
  assign _T_3168 = _T_2788 & _T_3167; // @[StoreQueue.scala 127:28:@1497.4]
  assign _T_3173 = _GEN_879 < 4'hd; // @[StoreQueue.scala 127:71:@1498.4]
  assign _T_3176 = _T_3173 & _T_2797; // @[StoreQueue.scala 127:79:@1500.4]
  assign _T_3178 = _T_3176 == 1'h0; // @[StoreQueue.scala 127:55:@1501.4]
  assign loadsToCheck_13 = _T_2861 ? _T_3168 : _T_3178; // @[StoreQueue.scala 126:83:@1502.4]
  assign _T_3190 = 4'he <= _GEN_879; // @[StoreQueue.scala 127:37:@1505.4]
  assign _T_3191 = _T_2805 & _T_3190; // @[StoreQueue.scala 127:28:@1506.4]
  assign _T_3196 = _GEN_879 < 4'he; // @[StoreQueue.scala 127:71:@1507.4]
  assign _T_3199 = _T_3196 & _T_2814; // @[StoreQueue.scala 127:79:@1509.4]
  assign _T_3201 = _T_3199 == 1'h0; // @[StoreQueue.scala 127:55:@1510.4]
  assign loadsToCheck_14 = _T_2861 ? _T_3191 : _T_3201; // @[StoreQueue.scala 126:83:@1511.4]
  assign _T_3213 = 4'hf <= _GEN_879; // @[StoreQueue.scala 127:37:@1514.4]
  assign loadsToCheck_15 = _T_2861 ? _T_3213 : 1'h1; // @[StoreQueue.scala 126:83:@1520.4]
  assign _T_3247 = loadsToCheck_0 & validEntriesInLoadQ_0; // @[StoreQueue.scala 133:16:@1538.4]
  assign _GEN_881 = 4'h1 == head ? checkBits_1 : checkBits_0; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_882 = 4'h2 == head ? checkBits_2 : _GEN_881; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_883 = 4'h3 == head ? checkBits_3 : _GEN_882; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_884 = 4'h4 == head ? checkBits_4 : _GEN_883; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_885 = 4'h5 == head ? checkBits_5 : _GEN_884; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_886 = 4'h6 == head ? checkBits_6 : _GEN_885; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_887 = 4'h7 == head ? checkBits_7 : _GEN_886; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_888 = 4'h8 == head ? checkBits_8 : _GEN_887; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_889 = 4'h9 == head ? checkBits_9 : _GEN_888; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_890 = 4'ha == head ? checkBits_10 : _GEN_889; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_891 = 4'hb == head ? checkBits_11 : _GEN_890; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_892 = 4'hc == head ? checkBits_12 : _GEN_891; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_893 = 4'hd == head ? checkBits_13 : _GEN_892; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_894 = 4'he == head ? checkBits_14 : _GEN_893; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_895 = 4'hf == head ? checkBits_15 : _GEN_894; // @[StoreQueue.scala 133:24:@1539.4]
  assign entriesToCheck_0 = _T_3247 & _GEN_895; // @[StoreQueue.scala 133:24:@1539.4]
  assign _T_3252 = loadsToCheck_1 & validEntriesInLoadQ_1; // @[StoreQueue.scala 133:16:@1540.4]
  assign entriesToCheck_1 = _T_3252 & _GEN_895; // @[StoreQueue.scala 133:24:@1541.4]
  assign _T_3257 = loadsToCheck_2 & validEntriesInLoadQ_2; // @[StoreQueue.scala 133:16:@1542.4]
  assign entriesToCheck_2 = _T_3257 & _GEN_895; // @[StoreQueue.scala 133:24:@1543.4]
  assign _T_3262 = loadsToCheck_3 & validEntriesInLoadQ_3; // @[StoreQueue.scala 133:16:@1544.4]
  assign entriesToCheck_3 = _T_3262 & _GEN_895; // @[StoreQueue.scala 133:24:@1545.4]
  assign _T_3267 = loadsToCheck_4 & validEntriesInLoadQ_4; // @[StoreQueue.scala 133:16:@1546.4]
  assign entriesToCheck_4 = _T_3267 & _GEN_895; // @[StoreQueue.scala 133:24:@1547.4]
  assign _T_3272 = loadsToCheck_5 & validEntriesInLoadQ_5; // @[StoreQueue.scala 133:16:@1548.4]
  assign entriesToCheck_5 = _T_3272 & _GEN_895; // @[StoreQueue.scala 133:24:@1549.4]
  assign _T_3277 = loadsToCheck_6 & validEntriesInLoadQ_6; // @[StoreQueue.scala 133:16:@1550.4]
  assign entriesToCheck_6 = _T_3277 & _GEN_895; // @[StoreQueue.scala 133:24:@1551.4]
  assign _T_3282 = loadsToCheck_7 & validEntriesInLoadQ_7; // @[StoreQueue.scala 133:16:@1552.4]
  assign entriesToCheck_7 = _T_3282 & _GEN_895; // @[StoreQueue.scala 133:24:@1553.4]
  assign _T_3287 = loadsToCheck_8 & validEntriesInLoadQ_8; // @[StoreQueue.scala 133:16:@1554.4]
  assign entriesToCheck_8 = _T_3287 & _GEN_895; // @[StoreQueue.scala 133:24:@1555.4]
  assign _T_3292 = loadsToCheck_9 & validEntriesInLoadQ_9; // @[StoreQueue.scala 133:16:@1556.4]
  assign entriesToCheck_9 = _T_3292 & _GEN_895; // @[StoreQueue.scala 133:24:@1557.4]
  assign _T_3297 = loadsToCheck_10 & validEntriesInLoadQ_10; // @[StoreQueue.scala 133:16:@1558.4]
  assign entriesToCheck_10 = _T_3297 & _GEN_895; // @[StoreQueue.scala 133:24:@1559.4]
  assign _T_3302 = loadsToCheck_11 & validEntriesInLoadQ_11; // @[StoreQueue.scala 133:16:@1560.4]
  assign entriesToCheck_11 = _T_3302 & _GEN_895; // @[StoreQueue.scala 133:24:@1561.4]
  assign _T_3307 = loadsToCheck_12 & validEntriesInLoadQ_12; // @[StoreQueue.scala 133:16:@1562.4]
  assign entriesToCheck_12 = _T_3307 & _GEN_895; // @[StoreQueue.scala 133:24:@1563.4]
  assign _T_3312 = loadsToCheck_13 & validEntriesInLoadQ_13; // @[StoreQueue.scala 133:16:@1564.4]
  assign entriesToCheck_13 = _T_3312 & _GEN_895; // @[StoreQueue.scala 133:24:@1565.4]
  assign _T_3317 = loadsToCheck_14 & validEntriesInLoadQ_14; // @[StoreQueue.scala 133:16:@1566.4]
  assign entriesToCheck_14 = _T_3317 & _GEN_895; // @[StoreQueue.scala 133:24:@1567.4]
  assign _T_3322 = loadsToCheck_15 & validEntriesInLoadQ_15; // @[StoreQueue.scala 133:16:@1568.4]
  assign entriesToCheck_15 = _T_3322 & _GEN_895; // @[StoreQueue.scala 133:24:@1569.4]
  assign _T_3370 = entriesToCheck_0 == 1'h0; // @[StoreQueue.scala 140:34:@1588.4]
  assign _T_3371 = _T_3370 | io_loadDataDone_0; // @[StoreQueue.scala 140:64:@1589.4]
  assign _GEN_897 = 4'h1 == head ? addrQ_1 : addrQ_0; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_898 = 4'h2 == head ? addrQ_2 : _GEN_897; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_899 = 4'h3 == head ? addrQ_3 : _GEN_898; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_900 = 4'h4 == head ? addrQ_4 : _GEN_899; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_901 = 4'h5 == head ? addrQ_5 : _GEN_900; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_902 = 4'h6 == head ? addrQ_6 : _GEN_901; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_903 = 4'h7 == head ? addrQ_7 : _GEN_902; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_904 = 4'h8 == head ? addrQ_8 : _GEN_903; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_905 = 4'h9 == head ? addrQ_9 : _GEN_904; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_906 = 4'ha == head ? addrQ_10 : _GEN_905; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_907 = 4'hb == head ? addrQ_11 : _GEN_906; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_908 = 4'hc == head ? addrQ_12 : _GEN_907; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_909 = 4'hd == head ? addrQ_13 : _GEN_908; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_910 = 4'he == head ? addrQ_14 : _GEN_909; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_911 = 4'hf == head ? addrQ_15 : _GEN_910; // @[StoreQueue.scala 141:51:@1590.4]
  assign _T_3375 = _GEN_911 != io_loadAddressQueue_0; // @[StoreQueue.scala 141:51:@1590.4]
  assign _T_3376 = io_loadAddressDone_0 & _T_3375; // @[StoreQueue.scala 141:36:@1591.4]
  assign noConflicts_0 = _T_3371 | _T_3376; // @[StoreQueue.scala 140:95:@1592.4]
  assign _T_3379 = entriesToCheck_1 == 1'h0; // @[StoreQueue.scala 140:34:@1594.4]
  assign _T_3380 = _T_3379 | io_loadDataDone_1; // @[StoreQueue.scala 140:64:@1595.4]
  assign _T_3384 = _GEN_911 != io_loadAddressQueue_1; // @[StoreQueue.scala 141:51:@1596.4]
  assign _T_3385 = io_loadAddressDone_1 & _T_3384; // @[StoreQueue.scala 141:36:@1597.4]
  assign noConflicts_1 = _T_3380 | _T_3385; // @[StoreQueue.scala 140:95:@1598.4]
  assign _T_3388 = entriesToCheck_2 == 1'h0; // @[StoreQueue.scala 140:34:@1600.4]
  assign _T_3389 = _T_3388 | io_loadDataDone_2; // @[StoreQueue.scala 140:64:@1601.4]
  assign _T_3393 = _GEN_911 != io_loadAddressQueue_2; // @[StoreQueue.scala 141:51:@1602.4]
  assign _T_3394 = io_loadAddressDone_2 & _T_3393; // @[StoreQueue.scala 141:36:@1603.4]
  assign noConflicts_2 = _T_3389 | _T_3394; // @[StoreQueue.scala 140:95:@1604.4]
  assign _T_3397 = entriesToCheck_3 == 1'h0; // @[StoreQueue.scala 140:34:@1606.4]
  assign _T_3398 = _T_3397 | io_loadDataDone_3; // @[StoreQueue.scala 140:64:@1607.4]
  assign _T_3402 = _GEN_911 != io_loadAddressQueue_3; // @[StoreQueue.scala 141:51:@1608.4]
  assign _T_3403 = io_loadAddressDone_3 & _T_3402; // @[StoreQueue.scala 141:36:@1609.4]
  assign noConflicts_3 = _T_3398 | _T_3403; // @[StoreQueue.scala 140:95:@1610.4]
  assign _T_3406 = entriesToCheck_4 == 1'h0; // @[StoreQueue.scala 140:34:@1612.4]
  assign _T_3407 = _T_3406 | io_loadDataDone_4; // @[StoreQueue.scala 140:64:@1613.4]
  assign _T_3411 = _GEN_911 != io_loadAddressQueue_4; // @[StoreQueue.scala 141:51:@1614.4]
  assign _T_3412 = io_loadAddressDone_4 & _T_3411; // @[StoreQueue.scala 141:36:@1615.4]
  assign noConflicts_4 = _T_3407 | _T_3412; // @[StoreQueue.scala 140:95:@1616.4]
  assign _T_3415 = entriesToCheck_5 == 1'h0; // @[StoreQueue.scala 140:34:@1618.4]
  assign _T_3416 = _T_3415 | io_loadDataDone_5; // @[StoreQueue.scala 140:64:@1619.4]
  assign _T_3420 = _GEN_911 != io_loadAddressQueue_5; // @[StoreQueue.scala 141:51:@1620.4]
  assign _T_3421 = io_loadAddressDone_5 & _T_3420; // @[StoreQueue.scala 141:36:@1621.4]
  assign noConflicts_5 = _T_3416 | _T_3421; // @[StoreQueue.scala 140:95:@1622.4]
  assign _T_3424 = entriesToCheck_6 == 1'h0; // @[StoreQueue.scala 140:34:@1624.4]
  assign _T_3425 = _T_3424 | io_loadDataDone_6; // @[StoreQueue.scala 140:64:@1625.4]
  assign _T_3429 = _GEN_911 != io_loadAddressQueue_6; // @[StoreQueue.scala 141:51:@1626.4]
  assign _T_3430 = io_loadAddressDone_6 & _T_3429; // @[StoreQueue.scala 141:36:@1627.4]
  assign noConflicts_6 = _T_3425 | _T_3430; // @[StoreQueue.scala 140:95:@1628.4]
  assign _T_3433 = entriesToCheck_7 == 1'h0; // @[StoreQueue.scala 140:34:@1630.4]
  assign _T_3434 = _T_3433 | io_loadDataDone_7; // @[StoreQueue.scala 140:64:@1631.4]
  assign _T_3438 = _GEN_911 != io_loadAddressQueue_7; // @[StoreQueue.scala 141:51:@1632.4]
  assign _T_3439 = io_loadAddressDone_7 & _T_3438; // @[StoreQueue.scala 141:36:@1633.4]
  assign noConflicts_7 = _T_3434 | _T_3439; // @[StoreQueue.scala 140:95:@1634.4]
  assign _T_3442 = entriesToCheck_8 == 1'h0; // @[StoreQueue.scala 140:34:@1636.4]
  assign _T_3443 = _T_3442 | io_loadDataDone_8; // @[StoreQueue.scala 140:64:@1637.4]
  assign _T_3447 = _GEN_911 != io_loadAddressQueue_8; // @[StoreQueue.scala 141:51:@1638.4]
  assign _T_3448 = io_loadAddressDone_8 & _T_3447; // @[StoreQueue.scala 141:36:@1639.4]
  assign noConflicts_8 = _T_3443 | _T_3448; // @[StoreQueue.scala 140:95:@1640.4]
  assign _T_3451 = entriesToCheck_9 == 1'h0; // @[StoreQueue.scala 140:34:@1642.4]
  assign _T_3452 = _T_3451 | io_loadDataDone_9; // @[StoreQueue.scala 140:64:@1643.4]
  assign _T_3456 = _GEN_911 != io_loadAddressQueue_9; // @[StoreQueue.scala 141:51:@1644.4]
  assign _T_3457 = io_loadAddressDone_9 & _T_3456; // @[StoreQueue.scala 141:36:@1645.4]
  assign noConflicts_9 = _T_3452 | _T_3457; // @[StoreQueue.scala 140:95:@1646.4]
  assign _T_3460 = entriesToCheck_10 == 1'h0; // @[StoreQueue.scala 140:34:@1648.4]
  assign _T_3461 = _T_3460 | io_loadDataDone_10; // @[StoreQueue.scala 140:64:@1649.4]
  assign _T_3465 = _GEN_911 != io_loadAddressQueue_10; // @[StoreQueue.scala 141:51:@1650.4]
  assign _T_3466 = io_loadAddressDone_10 & _T_3465; // @[StoreQueue.scala 141:36:@1651.4]
  assign noConflicts_10 = _T_3461 | _T_3466; // @[StoreQueue.scala 140:95:@1652.4]
  assign _T_3469 = entriesToCheck_11 == 1'h0; // @[StoreQueue.scala 140:34:@1654.4]
  assign _T_3470 = _T_3469 | io_loadDataDone_11; // @[StoreQueue.scala 140:64:@1655.4]
  assign _T_3474 = _GEN_911 != io_loadAddressQueue_11; // @[StoreQueue.scala 141:51:@1656.4]
  assign _T_3475 = io_loadAddressDone_11 & _T_3474; // @[StoreQueue.scala 141:36:@1657.4]
  assign noConflicts_11 = _T_3470 | _T_3475; // @[StoreQueue.scala 140:95:@1658.4]
  assign _T_3478 = entriesToCheck_12 == 1'h0; // @[StoreQueue.scala 140:34:@1660.4]
  assign _T_3479 = _T_3478 | io_loadDataDone_12; // @[StoreQueue.scala 140:64:@1661.4]
  assign _T_3483 = _GEN_911 != io_loadAddressQueue_12; // @[StoreQueue.scala 141:51:@1662.4]
  assign _T_3484 = io_loadAddressDone_12 & _T_3483; // @[StoreQueue.scala 141:36:@1663.4]
  assign noConflicts_12 = _T_3479 | _T_3484; // @[StoreQueue.scala 140:95:@1664.4]
  assign _T_3487 = entriesToCheck_13 == 1'h0; // @[StoreQueue.scala 140:34:@1666.4]
  assign _T_3488 = _T_3487 | io_loadDataDone_13; // @[StoreQueue.scala 140:64:@1667.4]
  assign _T_3492 = _GEN_911 != io_loadAddressQueue_13; // @[StoreQueue.scala 141:51:@1668.4]
  assign _T_3493 = io_loadAddressDone_13 & _T_3492; // @[StoreQueue.scala 141:36:@1669.4]
  assign noConflicts_13 = _T_3488 | _T_3493; // @[StoreQueue.scala 140:95:@1670.4]
  assign _T_3496 = entriesToCheck_14 == 1'h0; // @[StoreQueue.scala 140:34:@1672.4]
  assign _T_3497 = _T_3496 | io_loadDataDone_14; // @[StoreQueue.scala 140:64:@1673.4]
  assign _T_3501 = _GEN_911 != io_loadAddressQueue_14; // @[StoreQueue.scala 141:51:@1674.4]
  assign _T_3502 = io_loadAddressDone_14 & _T_3501; // @[StoreQueue.scala 141:36:@1675.4]
  assign noConflicts_14 = _T_3497 | _T_3502; // @[StoreQueue.scala 140:95:@1676.4]
  assign _T_3505 = entriesToCheck_15 == 1'h0; // @[StoreQueue.scala 140:34:@1678.4]
  assign _T_3506 = _T_3505 | io_loadDataDone_15; // @[StoreQueue.scala 140:64:@1679.4]
  assign _T_3510 = _GEN_911 != io_loadAddressQueue_15; // @[StoreQueue.scala 141:51:@1680.4]
  assign _T_3511 = io_loadAddressDone_15 & _T_3510; // @[StoreQueue.scala 141:36:@1681.4]
  assign noConflicts_15 = _T_3506 | _T_3511; // @[StoreQueue.scala 140:95:@1682.4]
  assign _GEN_913 = 4'h1 == head ? addrKnown_1 : addrKnown_0; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_914 = 4'h2 == head ? addrKnown_2 : _GEN_913; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_915 = 4'h3 == head ? addrKnown_3 : _GEN_914; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_916 = 4'h4 == head ? addrKnown_4 : _GEN_915; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_917 = 4'h5 == head ? addrKnown_5 : _GEN_916; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_918 = 4'h6 == head ? addrKnown_6 : _GEN_917; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_919 = 4'h7 == head ? addrKnown_7 : _GEN_918; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_920 = 4'h8 == head ? addrKnown_8 : _GEN_919; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_921 = 4'h9 == head ? addrKnown_9 : _GEN_920; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_922 = 4'ha == head ? addrKnown_10 : _GEN_921; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_923 = 4'hb == head ? addrKnown_11 : _GEN_922; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_924 = 4'hc == head ? addrKnown_12 : _GEN_923; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_925 = 4'hd == head ? addrKnown_13 : _GEN_924; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_926 = 4'he == head ? addrKnown_14 : _GEN_925; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_927 = 4'hf == head ? addrKnown_15 : _GEN_926; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_929 = 4'h1 == head ? dataKnown_1 : dataKnown_0; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_930 = 4'h2 == head ? dataKnown_2 : _GEN_929; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_931 = 4'h3 == head ? dataKnown_3 : _GEN_930; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_932 = 4'h4 == head ? dataKnown_4 : _GEN_931; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_933 = 4'h5 == head ? dataKnown_5 : _GEN_932; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_934 = 4'h6 == head ? dataKnown_6 : _GEN_933; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_935 = 4'h7 == head ? dataKnown_7 : _GEN_934; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_936 = 4'h8 == head ? dataKnown_8 : _GEN_935; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_937 = 4'h9 == head ? dataKnown_9 : _GEN_936; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_938 = 4'ha == head ? dataKnown_10 : _GEN_937; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_939 = 4'hb == head ? dataKnown_11 : _GEN_938; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_940 = 4'hc == head ? dataKnown_12 : _GEN_939; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_941 = 4'hd == head ? dataKnown_13 : _GEN_940; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_942 = 4'he == head ? dataKnown_14 : _GEN_941; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_943 = 4'hf == head ? dataKnown_15 : _GEN_942; // @[StoreQueue.scala 154:44:@1684.4]
  assign _T_3519 = _GEN_927 & _GEN_943; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_945 = 4'h1 == head ? storeCompleted_1 : storeCompleted_0; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_946 = 4'h2 == head ? storeCompleted_2 : _GEN_945; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_947 = 4'h3 == head ? storeCompleted_3 : _GEN_946; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_948 = 4'h4 == head ? storeCompleted_4 : _GEN_947; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_949 = 4'h5 == head ? storeCompleted_5 : _GEN_948; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_950 = 4'h6 == head ? storeCompleted_6 : _GEN_949; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_951 = 4'h7 == head ? storeCompleted_7 : _GEN_950; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_952 = 4'h8 == head ? storeCompleted_8 : _GEN_951; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_953 = 4'h9 == head ? storeCompleted_9 : _GEN_952; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_954 = 4'ha == head ? storeCompleted_10 : _GEN_953; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_955 = 4'hb == head ? storeCompleted_11 : _GEN_954; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_956 = 4'hc == head ? storeCompleted_12 : _GEN_955; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_957 = 4'hd == head ? storeCompleted_13 : _GEN_956; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_958 = 4'he == head ? storeCompleted_14 : _GEN_957; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_959 = 4'hf == head ? storeCompleted_15 : _GEN_958; // @[StoreQueue.scala 154:66:@1685.4]
  assign _T_3524 = _GEN_959 == 1'h0; // @[StoreQueue.scala 154:66:@1685.4]
  assign _T_3525 = _T_3519 & _T_3524; // @[StoreQueue.scala 154:63:@1686.4]
  assign _T_3528 = noConflicts_0 & noConflicts_1; // @[StoreQueue.scala 154:109:@1688.4]
  assign _T_3529 = _T_3528 & noConflicts_2; // @[StoreQueue.scala 154:109:@1689.4]
  assign _T_3530 = _T_3529 & noConflicts_3; // @[StoreQueue.scala 154:109:@1690.4]
  assign _T_3531 = _T_3530 & noConflicts_4; // @[StoreQueue.scala 154:109:@1691.4]
  assign _T_3532 = _T_3531 & noConflicts_5; // @[StoreQueue.scala 154:109:@1692.4]
  assign _T_3533 = _T_3532 & noConflicts_6; // @[StoreQueue.scala 154:109:@1693.4]
  assign _T_3534 = _T_3533 & noConflicts_7; // @[StoreQueue.scala 154:109:@1694.4]
  assign _T_3535 = _T_3534 & noConflicts_8; // @[StoreQueue.scala 154:109:@1695.4]
  assign _T_3536 = _T_3535 & noConflicts_9; // @[StoreQueue.scala 154:109:@1696.4]
  assign _T_3537 = _T_3536 & noConflicts_10; // @[StoreQueue.scala 154:109:@1697.4]
  assign _T_3538 = _T_3537 & noConflicts_11; // @[StoreQueue.scala 154:109:@1698.4]
  assign _T_3539 = _T_3538 & noConflicts_12; // @[StoreQueue.scala 154:109:@1699.4]
  assign _T_3540 = _T_3539 & noConflicts_13; // @[StoreQueue.scala 154:109:@1700.4]
  assign _T_3541 = _T_3540 & noConflicts_14; // @[StoreQueue.scala 154:109:@1701.4]
  assign _T_3542 = _T_3541 & noConflicts_15; // @[StoreQueue.scala 154:109:@1702.4]
  assign storeRequest = _T_3525 & _T_3542; // @[StoreQueue.scala 154:88:@1703.4]
  assign _T_3545 = head == 4'h0; // @[StoreQueue.scala 164:23:@1708.6]
  assign _T_3546 = _T_3545 & storeRequest; // @[StoreQueue.scala 164:43:@1709.6]
  assign _T_3547 = _T_3546 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1710.6]
  assign _GEN_960 = _T_3547 ? 1'h1 : storeCompleted_0; // @[StoreQueue.scala 164:86:@1711.6]
  assign _GEN_961 = initBits_0 ? 1'h0 : _GEN_960; // @[StoreQueue.scala 162:37:@1704.4]
  assign _T_3551 = head == 4'h1; // @[StoreQueue.scala 164:23:@1718.6]
  assign _T_3552 = _T_3551 & storeRequest; // @[StoreQueue.scala 164:43:@1719.6]
  assign _T_3553 = _T_3552 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1720.6]
  assign _GEN_962 = _T_3553 ? 1'h1 : storeCompleted_1; // @[StoreQueue.scala 164:86:@1721.6]
  assign _GEN_963 = initBits_1 ? 1'h0 : _GEN_962; // @[StoreQueue.scala 162:37:@1714.4]
  assign _T_3557 = head == 4'h2; // @[StoreQueue.scala 164:23:@1728.6]
  assign _T_3558 = _T_3557 & storeRequest; // @[StoreQueue.scala 164:43:@1729.6]
  assign _T_3559 = _T_3558 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1730.6]
  assign _GEN_964 = _T_3559 ? 1'h1 : storeCompleted_2; // @[StoreQueue.scala 164:86:@1731.6]
  assign _GEN_965 = initBits_2 ? 1'h0 : _GEN_964; // @[StoreQueue.scala 162:37:@1724.4]
  assign _T_3563 = head == 4'h3; // @[StoreQueue.scala 164:23:@1738.6]
  assign _T_3564 = _T_3563 & storeRequest; // @[StoreQueue.scala 164:43:@1739.6]
  assign _T_3565 = _T_3564 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1740.6]
  assign _GEN_966 = _T_3565 ? 1'h1 : storeCompleted_3; // @[StoreQueue.scala 164:86:@1741.6]
  assign _GEN_967 = initBits_3 ? 1'h0 : _GEN_966; // @[StoreQueue.scala 162:37:@1734.4]
  assign _T_3569 = head == 4'h4; // @[StoreQueue.scala 164:23:@1748.6]
  assign _T_3570 = _T_3569 & storeRequest; // @[StoreQueue.scala 164:43:@1749.6]
  assign _T_3571 = _T_3570 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1750.6]
  assign _GEN_968 = _T_3571 ? 1'h1 : storeCompleted_4; // @[StoreQueue.scala 164:86:@1751.6]
  assign _GEN_969 = initBits_4 ? 1'h0 : _GEN_968; // @[StoreQueue.scala 162:37:@1744.4]
  assign _T_3575 = head == 4'h5; // @[StoreQueue.scala 164:23:@1758.6]
  assign _T_3576 = _T_3575 & storeRequest; // @[StoreQueue.scala 164:43:@1759.6]
  assign _T_3577 = _T_3576 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1760.6]
  assign _GEN_970 = _T_3577 ? 1'h1 : storeCompleted_5; // @[StoreQueue.scala 164:86:@1761.6]
  assign _GEN_971 = initBits_5 ? 1'h0 : _GEN_970; // @[StoreQueue.scala 162:37:@1754.4]
  assign _T_3581 = head == 4'h6; // @[StoreQueue.scala 164:23:@1768.6]
  assign _T_3582 = _T_3581 & storeRequest; // @[StoreQueue.scala 164:43:@1769.6]
  assign _T_3583 = _T_3582 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1770.6]
  assign _GEN_972 = _T_3583 ? 1'h1 : storeCompleted_6; // @[StoreQueue.scala 164:86:@1771.6]
  assign _GEN_973 = initBits_6 ? 1'h0 : _GEN_972; // @[StoreQueue.scala 162:37:@1764.4]
  assign _T_3587 = head == 4'h7; // @[StoreQueue.scala 164:23:@1778.6]
  assign _T_3588 = _T_3587 & storeRequest; // @[StoreQueue.scala 164:43:@1779.6]
  assign _T_3589 = _T_3588 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1780.6]
  assign _GEN_974 = _T_3589 ? 1'h1 : storeCompleted_7; // @[StoreQueue.scala 164:86:@1781.6]
  assign _GEN_975 = initBits_7 ? 1'h0 : _GEN_974; // @[StoreQueue.scala 162:37:@1774.4]
  assign _T_3593 = head == 4'h8; // @[StoreQueue.scala 164:23:@1788.6]
  assign _T_3594 = _T_3593 & storeRequest; // @[StoreQueue.scala 164:43:@1789.6]
  assign _T_3595 = _T_3594 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1790.6]
  assign _GEN_976 = _T_3595 ? 1'h1 : storeCompleted_8; // @[StoreQueue.scala 164:86:@1791.6]
  assign _GEN_977 = initBits_8 ? 1'h0 : _GEN_976; // @[StoreQueue.scala 162:37:@1784.4]
  assign _T_3599 = head == 4'h9; // @[StoreQueue.scala 164:23:@1798.6]
  assign _T_3600 = _T_3599 & storeRequest; // @[StoreQueue.scala 164:43:@1799.6]
  assign _T_3601 = _T_3600 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1800.6]
  assign _GEN_978 = _T_3601 ? 1'h1 : storeCompleted_9; // @[StoreQueue.scala 164:86:@1801.6]
  assign _GEN_979 = initBits_9 ? 1'h0 : _GEN_978; // @[StoreQueue.scala 162:37:@1794.4]
  assign _T_3605 = head == 4'ha; // @[StoreQueue.scala 164:23:@1808.6]
  assign _T_3606 = _T_3605 & storeRequest; // @[StoreQueue.scala 164:43:@1809.6]
  assign _T_3607 = _T_3606 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1810.6]
  assign _GEN_980 = _T_3607 ? 1'h1 : storeCompleted_10; // @[StoreQueue.scala 164:86:@1811.6]
  assign _GEN_981 = initBits_10 ? 1'h0 : _GEN_980; // @[StoreQueue.scala 162:37:@1804.4]
  assign _T_3611 = head == 4'hb; // @[StoreQueue.scala 164:23:@1818.6]
  assign _T_3612 = _T_3611 & storeRequest; // @[StoreQueue.scala 164:43:@1819.6]
  assign _T_3613 = _T_3612 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1820.6]
  assign _GEN_982 = _T_3613 ? 1'h1 : storeCompleted_11; // @[StoreQueue.scala 164:86:@1821.6]
  assign _GEN_983 = initBits_11 ? 1'h0 : _GEN_982; // @[StoreQueue.scala 162:37:@1814.4]
  assign _T_3617 = head == 4'hc; // @[StoreQueue.scala 164:23:@1828.6]
  assign _T_3618 = _T_3617 & storeRequest; // @[StoreQueue.scala 164:43:@1829.6]
  assign _T_3619 = _T_3618 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1830.6]
  assign _GEN_984 = _T_3619 ? 1'h1 : storeCompleted_12; // @[StoreQueue.scala 164:86:@1831.6]
  assign _GEN_985 = initBits_12 ? 1'h0 : _GEN_984; // @[StoreQueue.scala 162:37:@1824.4]
  assign _T_3623 = head == 4'hd; // @[StoreQueue.scala 164:23:@1838.6]
  assign _T_3624 = _T_3623 & storeRequest; // @[StoreQueue.scala 164:43:@1839.6]
  assign _T_3625 = _T_3624 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1840.6]
  assign _GEN_986 = _T_3625 ? 1'h1 : storeCompleted_13; // @[StoreQueue.scala 164:86:@1841.6]
  assign _GEN_987 = initBits_13 ? 1'h0 : _GEN_986; // @[StoreQueue.scala 162:37:@1834.4]
  assign _T_3629 = head == 4'he; // @[StoreQueue.scala 164:23:@1848.6]
  assign _T_3630 = _T_3629 & storeRequest; // @[StoreQueue.scala 164:43:@1849.6]
  assign _T_3631 = _T_3630 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1850.6]
  assign _GEN_988 = _T_3631 ? 1'h1 : storeCompleted_14; // @[StoreQueue.scala 164:86:@1851.6]
  assign _GEN_989 = initBits_14 ? 1'h0 : _GEN_988; // @[StoreQueue.scala 162:37:@1844.4]
  assign _T_3635 = head == 4'hf; // @[StoreQueue.scala 164:23:@1858.6]
  assign _T_3636 = _T_3635 & storeRequest; // @[StoreQueue.scala 164:43:@1859.6]
  assign _T_3637 = _T_3636 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1860.6]
  assign _GEN_990 = _T_3637 ? 1'h1 : storeCompleted_15; // @[StoreQueue.scala 164:86:@1861.6]
  assign _GEN_991 = initBits_15 ? 1'h0 : _GEN_990; // @[StoreQueue.scala 162:37:@1854.4]
  assign entriesPorts_0_0 = portQ_0 == 1'h0; // @[StoreQueue.scala 180:72:@1865.4]
  assign entriesPorts_0_1 = portQ_1 == 1'h0; // @[StoreQueue.scala 180:72:@1867.4]
  assign entriesPorts_0_2 = portQ_2 == 1'h0; // @[StoreQueue.scala 180:72:@1869.4]
  assign entriesPorts_0_3 = portQ_3 == 1'h0; // @[StoreQueue.scala 180:72:@1871.4]
  assign entriesPorts_0_4 = portQ_4 == 1'h0; // @[StoreQueue.scala 180:72:@1873.4]
  assign entriesPorts_0_5 = portQ_5 == 1'h0; // @[StoreQueue.scala 180:72:@1875.4]
  assign entriesPorts_0_6 = portQ_6 == 1'h0; // @[StoreQueue.scala 180:72:@1877.4]
  assign entriesPorts_0_7 = portQ_7 == 1'h0; // @[StoreQueue.scala 180:72:@1879.4]
  assign entriesPorts_0_8 = portQ_8 == 1'h0; // @[StoreQueue.scala 180:72:@1881.4]
  assign entriesPorts_0_9 = portQ_9 == 1'h0; // @[StoreQueue.scala 180:72:@1883.4]
  assign entriesPorts_0_10 = portQ_10 == 1'h0; // @[StoreQueue.scala 180:72:@1885.4]
  assign entriesPorts_0_11 = portQ_11 == 1'h0; // @[StoreQueue.scala 180:72:@1887.4]
  assign entriesPorts_0_12 = portQ_12 == 1'h0; // @[StoreQueue.scala 180:72:@1889.4]
  assign entriesPorts_0_13 = portQ_13 == 1'h0; // @[StoreQueue.scala 180:72:@1891.4]
  assign entriesPorts_0_14 = portQ_14 == 1'h0; // @[StoreQueue.scala 180:72:@1893.4]
  assign entriesPorts_0_15 = portQ_15 == 1'h0; // @[StoreQueue.scala 180:72:@1895.4]
  assign _T_4122 = addrKnown_0 == 1'h0; // @[StoreQueue.scala 192:91:@1899.4]
  assign _T_4123 = entriesPorts_0_0 & _T_4122; // @[StoreQueue.scala 192:88:@1900.4]
  assign _T_4125 = addrKnown_1 == 1'h0; // @[StoreQueue.scala 192:91:@1901.4]
  assign _T_4126 = entriesPorts_0_1 & _T_4125; // @[StoreQueue.scala 192:88:@1902.4]
  assign _T_4128 = addrKnown_2 == 1'h0; // @[StoreQueue.scala 192:91:@1903.4]
  assign _T_4129 = entriesPorts_0_2 & _T_4128; // @[StoreQueue.scala 192:88:@1904.4]
  assign _T_4131 = addrKnown_3 == 1'h0; // @[StoreQueue.scala 192:91:@1905.4]
  assign _T_4132 = entriesPorts_0_3 & _T_4131; // @[StoreQueue.scala 192:88:@1906.4]
  assign _T_4134 = addrKnown_4 == 1'h0; // @[StoreQueue.scala 192:91:@1907.4]
  assign _T_4135 = entriesPorts_0_4 & _T_4134; // @[StoreQueue.scala 192:88:@1908.4]
  assign _T_4137 = addrKnown_5 == 1'h0; // @[StoreQueue.scala 192:91:@1909.4]
  assign _T_4138 = entriesPorts_0_5 & _T_4137; // @[StoreQueue.scala 192:88:@1910.4]
  assign _T_4140 = addrKnown_6 == 1'h0; // @[StoreQueue.scala 192:91:@1911.4]
  assign _T_4141 = entriesPorts_0_6 & _T_4140; // @[StoreQueue.scala 192:88:@1912.4]
  assign _T_4143 = addrKnown_7 == 1'h0; // @[StoreQueue.scala 192:91:@1913.4]
  assign _T_4144 = entriesPorts_0_7 & _T_4143; // @[StoreQueue.scala 192:88:@1914.4]
  assign _T_4146 = addrKnown_8 == 1'h0; // @[StoreQueue.scala 192:91:@1915.4]
  assign _T_4147 = entriesPorts_0_8 & _T_4146; // @[StoreQueue.scala 192:88:@1916.4]
  assign _T_4149 = addrKnown_9 == 1'h0; // @[StoreQueue.scala 192:91:@1917.4]
  assign _T_4150 = entriesPorts_0_9 & _T_4149; // @[StoreQueue.scala 192:88:@1918.4]
  assign _T_4152 = addrKnown_10 == 1'h0; // @[StoreQueue.scala 192:91:@1919.4]
  assign _T_4153 = entriesPorts_0_10 & _T_4152; // @[StoreQueue.scala 192:88:@1920.4]
  assign _T_4155 = addrKnown_11 == 1'h0; // @[StoreQueue.scala 192:91:@1921.4]
  assign _T_4156 = entriesPorts_0_11 & _T_4155; // @[StoreQueue.scala 192:88:@1922.4]
  assign _T_4158 = addrKnown_12 == 1'h0; // @[StoreQueue.scala 192:91:@1923.4]
  assign _T_4159 = entriesPorts_0_12 & _T_4158; // @[StoreQueue.scala 192:88:@1924.4]
  assign _T_4161 = addrKnown_13 == 1'h0; // @[StoreQueue.scala 192:91:@1925.4]
  assign _T_4162 = entriesPorts_0_13 & _T_4161; // @[StoreQueue.scala 192:88:@1926.4]
  assign _T_4164 = addrKnown_14 == 1'h0; // @[StoreQueue.scala 192:91:@1927.4]
  assign _T_4165 = entriesPorts_0_14 & _T_4164; // @[StoreQueue.scala 192:88:@1928.4]
  assign _T_4167 = addrKnown_15 == 1'h0; // @[StoreQueue.scala 192:91:@1929.4]
  assign _T_4168 = entriesPorts_0_15 & _T_4167; // @[StoreQueue.scala 192:88:@1930.4]
  assign _T_4192 = dataKnown_0 == 1'h0; // @[StoreQueue.scala 193:91:@1948.4]
  assign _T_4193 = entriesPorts_0_0 & _T_4192; // @[StoreQueue.scala 193:88:@1949.4]
  assign _T_4195 = dataKnown_1 == 1'h0; // @[StoreQueue.scala 193:91:@1950.4]
  assign _T_4196 = entriesPorts_0_1 & _T_4195; // @[StoreQueue.scala 193:88:@1951.4]
  assign _T_4198 = dataKnown_2 == 1'h0; // @[StoreQueue.scala 193:91:@1952.4]
  assign _T_4199 = entriesPorts_0_2 & _T_4198; // @[StoreQueue.scala 193:88:@1953.4]
  assign _T_4201 = dataKnown_3 == 1'h0; // @[StoreQueue.scala 193:91:@1954.4]
  assign _T_4202 = entriesPorts_0_3 & _T_4201; // @[StoreQueue.scala 193:88:@1955.4]
  assign _T_4204 = dataKnown_4 == 1'h0; // @[StoreQueue.scala 193:91:@1956.4]
  assign _T_4205 = entriesPorts_0_4 & _T_4204; // @[StoreQueue.scala 193:88:@1957.4]
  assign _T_4207 = dataKnown_5 == 1'h0; // @[StoreQueue.scala 193:91:@1958.4]
  assign _T_4208 = entriesPorts_0_5 & _T_4207; // @[StoreQueue.scala 193:88:@1959.4]
  assign _T_4210 = dataKnown_6 == 1'h0; // @[StoreQueue.scala 193:91:@1960.4]
  assign _T_4211 = entriesPorts_0_6 & _T_4210; // @[StoreQueue.scala 193:88:@1961.4]
  assign _T_4213 = dataKnown_7 == 1'h0; // @[StoreQueue.scala 193:91:@1962.4]
  assign _T_4214 = entriesPorts_0_7 & _T_4213; // @[StoreQueue.scala 193:88:@1963.4]
  assign _T_4216 = dataKnown_8 == 1'h0; // @[StoreQueue.scala 193:91:@1964.4]
  assign _T_4217 = entriesPorts_0_8 & _T_4216; // @[StoreQueue.scala 193:88:@1965.4]
  assign _T_4219 = dataKnown_9 == 1'h0; // @[StoreQueue.scala 193:91:@1966.4]
  assign _T_4220 = entriesPorts_0_9 & _T_4219; // @[StoreQueue.scala 193:88:@1967.4]
  assign _T_4222 = dataKnown_10 == 1'h0; // @[StoreQueue.scala 193:91:@1968.4]
  assign _T_4223 = entriesPorts_0_10 & _T_4222; // @[StoreQueue.scala 193:88:@1969.4]
  assign _T_4225 = dataKnown_11 == 1'h0; // @[StoreQueue.scala 193:91:@1970.4]
  assign _T_4226 = entriesPorts_0_11 & _T_4225; // @[StoreQueue.scala 193:88:@1971.4]
  assign _T_4228 = dataKnown_12 == 1'h0; // @[StoreQueue.scala 193:91:@1972.4]
  assign _T_4229 = entriesPorts_0_12 & _T_4228; // @[StoreQueue.scala 193:88:@1973.4]
  assign _T_4231 = dataKnown_13 == 1'h0; // @[StoreQueue.scala 193:91:@1974.4]
  assign _T_4232 = entriesPorts_0_13 & _T_4231; // @[StoreQueue.scala 193:88:@1975.4]
  assign _T_4234 = dataKnown_14 == 1'h0; // @[StoreQueue.scala 193:91:@1976.4]
  assign _T_4235 = entriesPorts_0_14 & _T_4234; // @[StoreQueue.scala 193:88:@1977.4]
  assign _T_4237 = dataKnown_15 == 1'h0; // @[StoreQueue.scala 193:91:@1978.4]
  assign _T_4238 = entriesPorts_0_15 & _T_4237; // @[StoreQueue.scala 193:88:@1979.4]
  assign _T_4263 = 16'h1 << head; // @[OneHot.scala 52:12:@1998.4]
  assign _T_4265 = _T_4263[0]; // @[util.scala 33:60:@2000.4]
  assign _T_4266 = _T_4263[1]; // @[util.scala 33:60:@2001.4]
  assign _T_4267 = _T_4263[2]; // @[util.scala 33:60:@2002.4]
  assign _T_4268 = _T_4263[3]; // @[util.scala 33:60:@2003.4]
  assign _T_4269 = _T_4263[4]; // @[util.scala 33:60:@2004.4]
  assign _T_4270 = _T_4263[5]; // @[util.scala 33:60:@2005.4]
  assign _T_4271 = _T_4263[6]; // @[util.scala 33:60:@2006.4]
  assign _T_4272 = _T_4263[7]; // @[util.scala 33:60:@2007.4]
  assign _T_4273 = _T_4263[8]; // @[util.scala 33:60:@2008.4]
  assign _T_4274 = _T_4263[9]; // @[util.scala 33:60:@2009.4]
  assign _T_4275 = _T_4263[10]; // @[util.scala 33:60:@2010.4]
  assign _T_4276 = _T_4263[11]; // @[util.scala 33:60:@2011.4]
  assign _T_4277 = _T_4263[12]; // @[util.scala 33:60:@2012.4]
  assign _T_4278 = _T_4263[13]; // @[util.scala 33:60:@2013.4]
  assign _T_4279 = _T_4263[14]; // @[util.scala 33:60:@2014.4]
  assign _T_4280 = _T_4263[15]; // @[util.scala 33:60:@2015.4]
  assign _T_4321 = _T_4168 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2033.4]
  assign _T_4322 = _T_4165 ? 16'h4000 : _T_4321; // @[Mux.scala 31:69:@2034.4]
  assign _T_4323 = _T_4162 ? 16'h2000 : _T_4322; // @[Mux.scala 31:69:@2035.4]
  assign _T_4324 = _T_4159 ? 16'h1000 : _T_4323; // @[Mux.scala 31:69:@2036.4]
  assign _T_4325 = _T_4156 ? 16'h800 : _T_4324; // @[Mux.scala 31:69:@2037.4]
  assign _T_4326 = _T_4153 ? 16'h400 : _T_4325; // @[Mux.scala 31:69:@2038.4]
  assign _T_4327 = _T_4150 ? 16'h200 : _T_4326; // @[Mux.scala 31:69:@2039.4]
  assign _T_4328 = _T_4147 ? 16'h100 : _T_4327; // @[Mux.scala 31:69:@2040.4]
  assign _T_4329 = _T_4144 ? 16'h80 : _T_4328; // @[Mux.scala 31:69:@2041.4]
  assign _T_4330 = _T_4141 ? 16'h40 : _T_4329; // @[Mux.scala 31:69:@2042.4]
  assign _T_4331 = _T_4138 ? 16'h20 : _T_4330; // @[Mux.scala 31:69:@2043.4]
  assign _T_4332 = _T_4135 ? 16'h10 : _T_4331; // @[Mux.scala 31:69:@2044.4]
  assign _T_4333 = _T_4132 ? 16'h8 : _T_4332; // @[Mux.scala 31:69:@2045.4]
  assign _T_4334 = _T_4129 ? 16'h4 : _T_4333; // @[Mux.scala 31:69:@2046.4]
  assign _T_4335 = _T_4126 ? 16'h2 : _T_4334; // @[Mux.scala 31:69:@2047.4]
  assign _T_4336 = _T_4123 ? 16'h1 : _T_4335; // @[Mux.scala 31:69:@2048.4]
  assign _T_4337 = _T_4336[0]; // @[OneHot.scala 66:30:@2049.4]
  assign _T_4338 = _T_4336[1]; // @[OneHot.scala 66:30:@2050.4]
  assign _T_4339 = _T_4336[2]; // @[OneHot.scala 66:30:@2051.4]
  assign _T_4340 = _T_4336[3]; // @[OneHot.scala 66:30:@2052.4]
  assign _T_4341 = _T_4336[4]; // @[OneHot.scala 66:30:@2053.4]
  assign _T_4342 = _T_4336[5]; // @[OneHot.scala 66:30:@2054.4]
  assign _T_4343 = _T_4336[6]; // @[OneHot.scala 66:30:@2055.4]
  assign _T_4344 = _T_4336[7]; // @[OneHot.scala 66:30:@2056.4]
  assign _T_4345 = _T_4336[8]; // @[OneHot.scala 66:30:@2057.4]
  assign _T_4346 = _T_4336[9]; // @[OneHot.scala 66:30:@2058.4]
  assign _T_4347 = _T_4336[10]; // @[OneHot.scala 66:30:@2059.4]
  assign _T_4348 = _T_4336[11]; // @[OneHot.scala 66:30:@2060.4]
  assign _T_4349 = _T_4336[12]; // @[OneHot.scala 66:30:@2061.4]
  assign _T_4350 = _T_4336[13]; // @[OneHot.scala 66:30:@2062.4]
  assign _T_4351 = _T_4336[14]; // @[OneHot.scala 66:30:@2063.4]
  assign _T_4352 = _T_4336[15]; // @[OneHot.scala 66:30:@2064.4]
  assign _T_4393 = _T_4123 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2082.4]
  assign _T_4394 = _T_4168 ? 16'h4000 : _T_4393; // @[Mux.scala 31:69:@2083.4]
  assign _T_4395 = _T_4165 ? 16'h2000 : _T_4394; // @[Mux.scala 31:69:@2084.4]
  assign _T_4396 = _T_4162 ? 16'h1000 : _T_4395; // @[Mux.scala 31:69:@2085.4]
  assign _T_4397 = _T_4159 ? 16'h800 : _T_4396; // @[Mux.scala 31:69:@2086.4]
  assign _T_4398 = _T_4156 ? 16'h400 : _T_4397; // @[Mux.scala 31:69:@2087.4]
  assign _T_4399 = _T_4153 ? 16'h200 : _T_4398; // @[Mux.scala 31:69:@2088.4]
  assign _T_4400 = _T_4150 ? 16'h100 : _T_4399; // @[Mux.scala 31:69:@2089.4]
  assign _T_4401 = _T_4147 ? 16'h80 : _T_4400; // @[Mux.scala 31:69:@2090.4]
  assign _T_4402 = _T_4144 ? 16'h40 : _T_4401; // @[Mux.scala 31:69:@2091.4]
  assign _T_4403 = _T_4141 ? 16'h20 : _T_4402; // @[Mux.scala 31:69:@2092.4]
  assign _T_4404 = _T_4138 ? 16'h10 : _T_4403; // @[Mux.scala 31:69:@2093.4]
  assign _T_4405 = _T_4135 ? 16'h8 : _T_4404; // @[Mux.scala 31:69:@2094.4]
  assign _T_4406 = _T_4132 ? 16'h4 : _T_4405; // @[Mux.scala 31:69:@2095.4]
  assign _T_4407 = _T_4129 ? 16'h2 : _T_4406; // @[Mux.scala 31:69:@2096.4]
  assign _T_4408 = _T_4126 ? 16'h1 : _T_4407; // @[Mux.scala 31:69:@2097.4]
  assign _T_4409 = _T_4408[0]; // @[OneHot.scala 66:30:@2098.4]
  assign _T_4410 = _T_4408[1]; // @[OneHot.scala 66:30:@2099.4]
  assign _T_4411 = _T_4408[2]; // @[OneHot.scala 66:30:@2100.4]
  assign _T_4412 = _T_4408[3]; // @[OneHot.scala 66:30:@2101.4]
  assign _T_4413 = _T_4408[4]; // @[OneHot.scala 66:30:@2102.4]
  assign _T_4414 = _T_4408[5]; // @[OneHot.scala 66:30:@2103.4]
  assign _T_4415 = _T_4408[6]; // @[OneHot.scala 66:30:@2104.4]
  assign _T_4416 = _T_4408[7]; // @[OneHot.scala 66:30:@2105.4]
  assign _T_4417 = _T_4408[8]; // @[OneHot.scala 66:30:@2106.4]
  assign _T_4418 = _T_4408[9]; // @[OneHot.scala 66:30:@2107.4]
  assign _T_4419 = _T_4408[10]; // @[OneHot.scala 66:30:@2108.4]
  assign _T_4420 = _T_4408[11]; // @[OneHot.scala 66:30:@2109.4]
  assign _T_4421 = _T_4408[12]; // @[OneHot.scala 66:30:@2110.4]
  assign _T_4422 = _T_4408[13]; // @[OneHot.scala 66:30:@2111.4]
  assign _T_4423 = _T_4408[14]; // @[OneHot.scala 66:30:@2112.4]
  assign _T_4424 = _T_4408[15]; // @[OneHot.scala 66:30:@2113.4]
  assign _T_4465 = _T_4126 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2131.4]
  assign _T_4466 = _T_4123 ? 16'h4000 : _T_4465; // @[Mux.scala 31:69:@2132.4]
  assign _T_4467 = _T_4168 ? 16'h2000 : _T_4466; // @[Mux.scala 31:69:@2133.4]
  assign _T_4468 = _T_4165 ? 16'h1000 : _T_4467; // @[Mux.scala 31:69:@2134.4]
  assign _T_4469 = _T_4162 ? 16'h800 : _T_4468; // @[Mux.scala 31:69:@2135.4]
  assign _T_4470 = _T_4159 ? 16'h400 : _T_4469; // @[Mux.scala 31:69:@2136.4]
  assign _T_4471 = _T_4156 ? 16'h200 : _T_4470; // @[Mux.scala 31:69:@2137.4]
  assign _T_4472 = _T_4153 ? 16'h100 : _T_4471; // @[Mux.scala 31:69:@2138.4]
  assign _T_4473 = _T_4150 ? 16'h80 : _T_4472; // @[Mux.scala 31:69:@2139.4]
  assign _T_4474 = _T_4147 ? 16'h40 : _T_4473; // @[Mux.scala 31:69:@2140.4]
  assign _T_4475 = _T_4144 ? 16'h20 : _T_4474; // @[Mux.scala 31:69:@2141.4]
  assign _T_4476 = _T_4141 ? 16'h10 : _T_4475; // @[Mux.scala 31:69:@2142.4]
  assign _T_4477 = _T_4138 ? 16'h8 : _T_4476; // @[Mux.scala 31:69:@2143.4]
  assign _T_4478 = _T_4135 ? 16'h4 : _T_4477; // @[Mux.scala 31:69:@2144.4]
  assign _T_4479 = _T_4132 ? 16'h2 : _T_4478; // @[Mux.scala 31:69:@2145.4]
  assign _T_4480 = _T_4129 ? 16'h1 : _T_4479; // @[Mux.scala 31:69:@2146.4]
  assign _T_4481 = _T_4480[0]; // @[OneHot.scala 66:30:@2147.4]
  assign _T_4482 = _T_4480[1]; // @[OneHot.scala 66:30:@2148.4]
  assign _T_4483 = _T_4480[2]; // @[OneHot.scala 66:30:@2149.4]
  assign _T_4484 = _T_4480[3]; // @[OneHot.scala 66:30:@2150.4]
  assign _T_4485 = _T_4480[4]; // @[OneHot.scala 66:30:@2151.4]
  assign _T_4486 = _T_4480[5]; // @[OneHot.scala 66:30:@2152.4]
  assign _T_4487 = _T_4480[6]; // @[OneHot.scala 66:30:@2153.4]
  assign _T_4488 = _T_4480[7]; // @[OneHot.scala 66:30:@2154.4]
  assign _T_4489 = _T_4480[8]; // @[OneHot.scala 66:30:@2155.4]
  assign _T_4490 = _T_4480[9]; // @[OneHot.scala 66:30:@2156.4]
  assign _T_4491 = _T_4480[10]; // @[OneHot.scala 66:30:@2157.4]
  assign _T_4492 = _T_4480[11]; // @[OneHot.scala 66:30:@2158.4]
  assign _T_4493 = _T_4480[12]; // @[OneHot.scala 66:30:@2159.4]
  assign _T_4494 = _T_4480[13]; // @[OneHot.scala 66:30:@2160.4]
  assign _T_4495 = _T_4480[14]; // @[OneHot.scala 66:30:@2161.4]
  assign _T_4496 = _T_4480[15]; // @[OneHot.scala 66:30:@2162.4]
  assign _T_4537 = _T_4129 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2180.4]
  assign _T_4538 = _T_4126 ? 16'h4000 : _T_4537; // @[Mux.scala 31:69:@2181.4]
  assign _T_4539 = _T_4123 ? 16'h2000 : _T_4538; // @[Mux.scala 31:69:@2182.4]
  assign _T_4540 = _T_4168 ? 16'h1000 : _T_4539; // @[Mux.scala 31:69:@2183.4]
  assign _T_4541 = _T_4165 ? 16'h800 : _T_4540; // @[Mux.scala 31:69:@2184.4]
  assign _T_4542 = _T_4162 ? 16'h400 : _T_4541; // @[Mux.scala 31:69:@2185.4]
  assign _T_4543 = _T_4159 ? 16'h200 : _T_4542; // @[Mux.scala 31:69:@2186.4]
  assign _T_4544 = _T_4156 ? 16'h100 : _T_4543; // @[Mux.scala 31:69:@2187.4]
  assign _T_4545 = _T_4153 ? 16'h80 : _T_4544; // @[Mux.scala 31:69:@2188.4]
  assign _T_4546 = _T_4150 ? 16'h40 : _T_4545; // @[Mux.scala 31:69:@2189.4]
  assign _T_4547 = _T_4147 ? 16'h20 : _T_4546; // @[Mux.scala 31:69:@2190.4]
  assign _T_4548 = _T_4144 ? 16'h10 : _T_4547; // @[Mux.scala 31:69:@2191.4]
  assign _T_4549 = _T_4141 ? 16'h8 : _T_4548; // @[Mux.scala 31:69:@2192.4]
  assign _T_4550 = _T_4138 ? 16'h4 : _T_4549; // @[Mux.scala 31:69:@2193.4]
  assign _T_4551 = _T_4135 ? 16'h2 : _T_4550; // @[Mux.scala 31:69:@2194.4]
  assign _T_4552 = _T_4132 ? 16'h1 : _T_4551; // @[Mux.scala 31:69:@2195.4]
  assign _T_4553 = _T_4552[0]; // @[OneHot.scala 66:30:@2196.4]
  assign _T_4554 = _T_4552[1]; // @[OneHot.scala 66:30:@2197.4]
  assign _T_4555 = _T_4552[2]; // @[OneHot.scala 66:30:@2198.4]
  assign _T_4556 = _T_4552[3]; // @[OneHot.scala 66:30:@2199.4]
  assign _T_4557 = _T_4552[4]; // @[OneHot.scala 66:30:@2200.4]
  assign _T_4558 = _T_4552[5]; // @[OneHot.scala 66:30:@2201.4]
  assign _T_4559 = _T_4552[6]; // @[OneHot.scala 66:30:@2202.4]
  assign _T_4560 = _T_4552[7]; // @[OneHot.scala 66:30:@2203.4]
  assign _T_4561 = _T_4552[8]; // @[OneHot.scala 66:30:@2204.4]
  assign _T_4562 = _T_4552[9]; // @[OneHot.scala 66:30:@2205.4]
  assign _T_4563 = _T_4552[10]; // @[OneHot.scala 66:30:@2206.4]
  assign _T_4564 = _T_4552[11]; // @[OneHot.scala 66:30:@2207.4]
  assign _T_4565 = _T_4552[12]; // @[OneHot.scala 66:30:@2208.4]
  assign _T_4566 = _T_4552[13]; // @[OneHot.scala 66:30:@2209.4]
  assign _T_4567 = _T_4552[14]; // @[OneHot.scala 66:30:@2210.4]
  assign _T_4568 = _T_4552[15]; // @[OneHot.scala 66:30:@2211.4]
  assign _T_4609 = _T_4132 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2229.4]
  assign _T_4610 = _T_4129 ? 16'h4000 : _T_4609; // @[Mux.scala 31:69:@2230.4]
  assign _T_4611 = _T_4126 ? 16'h2000 : _T_4610; // @[Mux.scala 31:69:@2231.4]
  assign _T_4612 = _T_4123 ? 16'h1000 : _T_4611; // @[Mux.scala 31:69:@2232.4]
  assign _T_4613 = _T_4168 ? 16'h800 : _T_4612; // @[Mux.scala 31:69:@2233.4]
  assign _T_4614 = _T_4165 ? 16'h400 : _T_4613; // @[Mux.scala 31:69:@2234.4]
  assign _T_4615 = _T_4162 ? 16'h200 : _T_4614; // @[Mux.scala 31:69:@2235.4]
  assign _T_4616 = _T_4159 ? 16'h100 : _T_4615; // @[Mux.scala 31:69:@2236.4]
  assign _T_4617 = _T_4156 ? 16'h80 : _T_4616; // @[Mux.scala 31:69:@2237.4]
  assign _T_4618 = _T_4153 ? 16'h40 : _T_4617; // @[Mux.scala 31:69:@2238.4]
  assign _T_4619 = _T_4150 ? 16'h20 : _T_4618; // @[Mux.scala 31:69:@2239.4]
  assign _T_4620 = _T_4147 ? 16'h10 : _T_4619; // @[Mux.scala 31:69:@2240.4]
  assign _T_4621 = _T_4144 ? 16'h8 : _T_4620; // @[Mux.scala 31:69:@2241.4]
  assign _T_4622 = _T_4141 ? 16'h4 : _T_4621; // @[Mux.scala 31:69:@2242.4]
  assign _T_4623 = _T_4138 ? 16'h2 : _T_4622; // @[Mux.scala 31:69:@2243.4]
  assign _T_4624 = _T_4135 ? 16'h1 : _T_4623; // @[Mux.scala 31:69:@2244.4]
  assign _T_4625 = _T_4624[0]; // @[OneHot.scala 66:30:@2245.4]
  assign _T_4626 = _T_4624[1]; // @[OneHot.scala 66:30:@2246.4]
  assign _T_4627 = _T_4624[2]; // @[OneHot.scala 66:30:@2247.4]
  assign _T_4628 = _T_4624[3]; // @[OneHot.scala 66:30:@2248.4]
  assign _T_4629 = _T_4624[4]; // @[OneHot.scala 66:30:@2249.4]
  assign _T_4630 = _T_4624[5]; // @[OneHot.scala 66:30:@2250.4]
  assign _T_4631 = _T_4624[6]; // @[OneHot.scala 66:30:@2251.4]
  assign _T_4632 = _T_4624[7]; // @[OneHot.scala 66:30:@2252.4]
  assign _T_4633 = _T_4624[8]; // @[OneHot.scala 66:30:@2253.4]
  assign _T_4634 = _T_4624[9]; // @[OneHot.scala 66:30:@2254.4]
  assign _T_4635 = _T_4624[10]; // @[OneHot.scala 66:30:@2255.4]
  assign _T_4636 = _T_4624[11]; // @[OneHot.scala 66:30:@2256.4]
  assign _T_4637 = _T_4624[12]; // @[OneHot.scala 66:30:@2257.4]
  assign _T_4638 = _T_4624[13]; // @[OneHot.scala 66:30:@2258.4]
  assign _T_4639 = _T_4624[14]; // @[OneHot.scala 66:30:@2259.4]
  assign _T_4640 = _T_4624[15]; // @[OneHot.scala 66:30:@2260.4]
  assign _T_4681 = _T_4135 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2278.4]
  assign _T_4682 = _T_4132 ? 16'h4000 : _T_4681; // @[Mux.scala 31:69:@2279.4]
  assign _T_4683 = _T_4129 ? 16'h2000 : _T_4682; // @[Mux.scala 31:69:@2280.4]
  assign _T_4684 = _T_4126 ? 16'h1000 : _T_4683; // @[Mux.scala 31:69:@2281.4]
  assign _T_4685 = _T_4123 ? 16'h800 : _T_4684; // @[Mux.scala 31:69:@2282.4]
  assign _T_4686 = _T_4168 ? 16'h400 : _T_4685; // @[Mux.scala 31:69:@2283.4]
  assign _T_4687 = _T_4165 ? 16'h200 : _T_4686; // @[Mux.scala 31:69:@2284.4]
  assign _T_4688 = _T_4162 ? 16'h100 : _T_4687; // @[Mux.scala 31:69:@2285.4]
  assign _T_4689 = _T_4159 ? 16'h80 : _T_4688; // @[Mux.scala 31:69:@2286.4]
  assign _T_4690 = _T_4156 ? 16'h40 : _T_4689; // @[Mux.scala 31:69:@2287.4]
  assign _T_4691 = _T_4153 ? 16'h20 : _T_4690; // @[Mux.scala 31:69:@2288.4]
  assign _T_4692 = _T_4150 ? 16'h10 : _T_4691; // @[Mux.scala 31:69:@2289.4]
  assign _T_4693 = _T_4147 ? 16'h8 : _T_4692; // @[Mux.scala 31:69:@2290.4]
  assign _T_4694 = _T_4144 ? 16'h4 : _T_4693; // @[Mux.scala 31:69:@2291.4]
  assign _T_4695 = _T_4141 ? 16'h2 : _T_4694; // @[Mux.scala 31:69:@2292.4]
  assign _T_4696 = _T_4138 ? 16'h1 : _T_4695; // @[Mux.scala 31:69:@2293.4]
  assign _T_4697 = _T_4696[0]; // @[OneHot.scala 66:30:@2294.4]
  assign _T_4698 = _T_4696[1]; // @[OneHot.scala 66:30:@2295.4]
  assign _T_4699 = _T_4696[2]; // @[OneHot.scala 66:30:@2296.4]
  assign _T_4700 = _T_4696[3]; // @[OneHot.scala 66:30:@2297.4]
  assign _T_4701 = _T_4696[4]; // @[OneHot.scala 66:30:@2298.4]
  assign _T_4702 = _T_4696[5]; // @[OneHot.scala 66:30:@2299.4]
  assign _T_4703 = _T_4696[6]; // @[OneHot.scala 66:30:@2300.4]
  assign _T_4704 = _T_4696[7]; // @[OneHot.scala 66:30:@2301.4]
  assign _T_4705 = _T_4696[8]; // @[OneHot.scala 66:30:@2302.4]
  assign _T_4706 = _T_4696[9]; // @[OneHot.scala 66:30:@2303.4]
  assign _T_4707 = _T_4696[10]; // @[OneHot.scala 66:30:@2304.4]
  assign _T_4708 = _T_4696[11]; // @[OneHot.scala 66:30:@2305.4]
  assign _T_4709 = _T_4696[12]; // @[OneHot.scala 66:30:@2306.4]
  assign _T_4710 = _T_4696[13]; // @[OneHot.scala 66:30:@2307.4]
  assign _T_4711 = _T_4696[14]; // @[OneHot.scala 66:30:@2308.4]
  assign _T_4712 = _T_4696[15]; // @[OneHot.scala 66:30:@2309.4]
  assign _T_4753 = _T_4138 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2327.4]
  assign _T_4754 = _T_4135 ? 16'h4000 : _T_4753; // @[Mux.scala 31:69:@2328.4]
  assign _T_4755 = _T_4132 ? 16'h2000 : _T_4754; // @[Mux.scala 31:69:@2329.4]
  assign _T_4756 = _T_4129 ? 16'h1000 : _T_4755; // @[Mux.scala 31:69:@2330.4]
  assign _T_4757 = _T_4126 ? 16'h800 : _T_4756; // @[Mux.scala 31:69:@2331.4]
  assign _T_4758 = _T_4123 ? 16'h400 : _T_4757; // @[Mux.scala 31:69:@2332.4]
  assign _T_4759 = _T_4168 ? 16'h200 : _T_4758; // @[Mux.scala 31:69:@2333.4]
  assign _T_4760 = _T_4165 ? 16'h100 : _T_4759; // @[Mux.scala 31:69:@2334.4]
  assign _T_4761 = _T_4162 ? 16'h80 : _T_4760; // @[Mux.scala 31:69:@2335.4]
  assign _T_4762 = _T_4159 ? 16'h40 : _T_4761; // @[Mux.scala 31:69:@2336.4]
  assign _T_4763 = _T_4156 ? 16'h20 : _T_4762; // @[Mux.scala 31:69:@2337.4]
  assign _T_4764 = _T_4153 ? 16'h10 : _T_4763; // @[Mux.scala 31:69:@2338.4]
  assign _T_4765 = _T_4150 ? 16'h8 : _T_4764; // @[Mux.scala 31:69:@2339.4]
  assign _T_4766 = _T_4147 ? 16'h4 : _T_4765; // @[Mux.scala 31:69:@2340.4]
  assign _T_4767 = _T_4144 ? 16'h2 : _T_4766; // @[Mux.scala 31:69:@2341.4]
  assign _T_4768 = _T_4141 ? 16'h1 : _T_4767; // @[Mux.scala 31:69:@2342.4]
  assign _T_4769 = _T_4768[0]; // @[OneHot.scala 66:30:@2343.4]
  assign _T_4770 = _T_4768[1]; // @[OneHot.scala 66:30:@2344.4]
  assign _T_4771 = _T_4768[2]; // @[OneHot.scala 66:30:@2345.4]
  assign _T_4772 = _T_4768[3]; // @[OneHot.scala 66:30:@2346.4]
  assign _T_4773 = _T_4768[4]; // @[OneHot.scala 66:30:@2347.4]
  assign _T_4774 = _T_4768[5]; // @[OneHot.scala 66:30:@2348.4]
  assign _T_4775 = _T_4768[6]; // @[OneHot.scala 66:30:@2349.4]
  assign _T_4776 = _T_4768[7]; // @[OneHot.scala 66:30:@2350.4]
  assign _T_4777 = _T_4768[8]; // @[OneHot.scala 66:30:@2351.4]
  assign _T_4778 = _T_4768[9]; // @[OneHot.scala 66:30:@2352.4]
  assign _T_4779 = _T_4768[10]; // @[OneHot.scala 66:30:@2353.4]
  assign _T_4780 = _T_4768[11]; // @[OneHot.scala 66:30:@2354.4]
  assign _T_4781 = _T_4768[12]; // @[OneHot.scala 66:30:@2355.4]
  assign _T_4782 = _T_4768[13]; // @[OneHot.scala 66:30:@2356.4]
  assign _T_4783 = _T_4768[14]; // @[OneHot.scala 66:30:@2357.4]
  assign _T_4784 = _T_4768[15]; // @[OneHot.scala 66:30:@2358.4]
  assign _T_4825 = _T_4141 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2376.4]
  assign _T_4826 = _T_4138 ? 16'h4000 : _T_4825; // @[Mux.scala 31:69:@2377.4]
  assign _T_4827 = _T_4135 ? 16'h2000 : _T_4826; // @[Mux.scala 31:69:@2378.4]
  assign _T_4828 = _T_4132 ? 16'h1000 : _T_4827; // @[Mux.scala 31:69:@2379.4]
  assign _T_4829 = _T_4129 ? 16'h800 : _T_4828; // @[Mux.scala 31:69:@2380.4]
  assign _T_4830 = _T_4126 ? 16'h400 : _T_4829; // @[Mux.scala 31:69:@2381.4]
  assign _T_4831 = _T_4123 ? 16'h200 : _T_4830; // @[Mux.scala 31:69:@2382.4]
  assign _T_4832 = _T_4168 ? 16'h100 : _T_4831; // @[Mux.scala 31:69:@2383.4]
  assign _T_4833 = _T_4165 ? 16'h80 : _T_4832; // @[Mux.scala 31:69:@2384.4]
  assign _T_4834 = _T_4162 ? 16'h40 : _T_4833; // @[Mux.scala 31:69:@2385.4]
  assign _T_4835 = _T_4159 ? 16'h20 : _T_4834; // @[Mux.scala 31:69:@2386.4]
  assign _T_4836 = _T_4156 ? 16'h10 : _T_4835; // @[Mux.scala 31:69:@2387.4]
  assign _T_4837 = _T_4153 ? 16'h8 : _T_4836; // @[Mux.scala 31:69:@2388.4]
  assign _T_4838 = _T_4150 ? 16'h4 : _T_4837; // @[Mux.scala 31:69:@2389.4]
  assign _T_4839 = _T_4147 ? 16'h2 : _T_4838; // @[Mux.scala 31:69:@2390.4]
  assign _T_4840 = _T_4144 ? 16'h1 : _T_4839; // @[Mux.scala 31:69:@2391.4]
  assign _T_4841 = _T_4840[0]; // @[OneHot.scala 66:30:@2392.4]
  assign _T_4842 = _T_4840[1]; // @[OneHot.scala 66:30:@2393.4]
  assign _T_4843 = _T_4840[2]; // @[OneHot.scala 66:30:@2394.4]
  assign _T_4844 = _T_4840[3]; // @[OneHot.scala 66:30:@2395.4]
  assign _T_4845 = _T_4840[4]; // @[OneHot.scala 66:30:@2396.4]
  assign _T_4846 = _T_4840[5]; // @[OneHot.scala 66:30:@2397.4]
  assign _T_4847 = _T_4840[6]; // @[OneHot.scala 66:30:@2398.4]
  assign _T_4848 = _T_4840[7]; // @[OneHot.scala 66:30:@2399.4]
  assign _T_4849 = _T_4840[8]; // @[OneHot.scala 66:30:@2400.4]
  assign _T_4850 = _T_4840[9]; // @[OneHot.scala 66:30:@2401.4]
  assign _T_4851 = _T_4840[10]; // @[OneHot.scala 66:30:@2402.4]
  assign _T_4852 = _T_4840[11]; // @[OneHot.scala 66:30:@2403.4]
  assign _T_4853 = _T_4840[12]; // @[OneHot.scala 66:30:@2404.4]
  assign _T_4854 = _T_4840[13]; // @[OneHot.scala 66:30:@2405.4]
  assign _T_4855 = _T_4840[14]; // @[OneHot.scala 66:30:@2406.4]
  assign _T_4856 = _T_4840[15]; // @[OneHot.scala 66:30:@2407.4]
  assign _T_4897 = _T_4144 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2425.4]
  assign _T_4898 = _T_4141 ? 16'h4000 : _T_4897; // @[Mux.scala 31:69:@2426.4]
  assign _T_4899 = _T_4138 ? 16'h2000 : _T_4898; // @[Mux.scala 31:69:@2427.4]
  assign _T_4900 = _T_4135 ? 16'h1000 : _T_4899; // @[Mux.scala 31:69:@2428.4]
  assign _T_4901 = _T_4132 ? 16'h800 : _T_4900; // @[Mux.scala 31:69:@2429.4]
  assign _T_4902 = _T_4129 ? 16'h400 : _T_4901; // @[Mux.scala 31:69:@2430.4]
  assign _T_4903 = _T_4126 ? 16'h200 : _T_4902; // @[Mux.scala 31:69:@2431.4]
  assign _T_4904 = _T_4123 ? 16'h100 : _T_4903; // @[Mux.scala 31:69:@2432.4]
  assign _T_4905 = _T_4168 ? 16'h80 : _T_4904; // @[Mux.scala 31:69:@2433.4]
  assign _T_4906 = _T_4165 ? 16'h40 : _T_4905; // @[Mux.scala 31:69:@2434.4]
  assign _T_4907 = _T_4162 ? 16'h20 : _T_4906; // @[Mux.scala 31:69:@2435.4]
  assign _T_4908 = _T_4159 ? 16'h10 : _T_4907; // @[Mux.scala 31:69:@2436.4]
  assign _T_4909 = _T_4156 ? 16'h8 : _T_4908; // @[Mux.scala 31:69:@2437.4]
  assign _T_4910 = _T_4153 ? 16'h4 : _T_4909; // @[Mux.scala 31:69:@2438.4]
  assign _T_4911 = _T_4150 ? 16'h2 : _T_4910; // @[Mux.scala 31:69:@2439.4]
  assign _T_4912 = _T_4147 ? 16'h1 : _T_4911; // @[Mux.scala 31:69:@2440.4]
  assign _T_4913 = _T_4912[0]; // @[OneHot.scala 66:30:@2441.4]
  assign _T_4914 = _T_4912[1]; // @[OneHot.scala 66:30:@2442.4]
  assign _T_4915 = _T_4912[2]; // @[OneHot.scala 66:30:@2443.4]
  assign _T_4916 = _T_4912[3]; // @[OneHot.scala 66:30:@2444.4]
  assign _T_4917 = _T_4912[4]; // @[OneHot.scala 66:30:@2445.4]
  assign _T_4918 = _T_4912[5]; // @[OneHot.scala 66:30:@2446.4]
  assign _T_4919 = _T_4912[6]; // @[OneHot.scala 66:30:@2447.4]
  assign _T_4920 = _T_4912[7]; // @[OneHot.scala 66:30:@2448.4]
  assign _T_4921 = _T_4912[8]; // @[OneHot.scala 66:30:@2449.4]
  assign _T_4922 = _T_4912[9]; // @[OneHot.scala 66:30:@2450.4]
  assign _T_4923 = _T_4912[10]; // @[OneHot.scala 66:30:@2451.4]
  assign _T_4924 = _T_4912[11]; // @[OneHot.scala 66:30:@2452.4]
  assign _T_4925 = _T_4912[12]; // @[OneHot.scala 66:30:@2453.4]
  assign _T_4926 = _T_4912[13]; // @[OneHot.scala 66:30:@2454.4]
  assign _T_4927 = _T_4912[14]; // @[OneHot.scala 66:30:@2455.4]
  assign _T_4928 = _T_4912[15]; // @[OneHot.scala 66:30:@2456.4]
  assign _T_4969 = _T_4147 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2474.4]
  assign _T_4970 = _T_4144 ? 16'h4000 : _T_4969; // @[Mux.scala 31:69:@2475.4]
  assign _T_4971 = _T_4141 ? 16'h2000 : _T_4970; // @[Mux.scala 31:69:@2476.4]
  assign _T_4972 = _T_4138 ? 16'h1000 : _T_4971; // @[Mux.scala 31:69:@2477.4]
  assign _T_4973 = _T_4135 ? 16'h800 : _T_4972; // @[Mux.scala 31:69:@2478.4]
  assign _T_4974 = _T_4132 ? 16'h400 : _T_4973; // @[Mux.scala 31:69:@2479.4]
  assign _T_4975 = _T_4129 ? 16'h200 : _T_4974; // @[Mux.scala 31:69:@2480.4]
  assign _T_4976 = _T_4126 ? 16'h100 : _T_4975; // @[Mux.scala 31:69:@2481.4]
  assign _T_4977 = _T_4123 ? 16'h80 : _T_4976; // @[Mux.scala 31:69:@2482.4]
  assign _T_4978 = _T_4168 ? 16'h40 : _T_4977; // @[Mux.scala 31:69:@2483.4]
  assign _T_4979 = _T_4165 ? 16'h20 : _T_4978; // @[Mux.scala 31:69:@2484.4]
  assign _T_4980 = _T_4162 ? 16'h10 : _T_4979; // @[Mux.scala 31:69:@2485.4]
  assign _T_4981 = _T_4159 ? 16'h8 : _T_4980; // @[Mux.scala 31:69:@2486.4]
  assign _T_4982 = _T_4156 ? 16'h4 : _T_4981; // @[Mux.scala 31:69:@2487.4]
  assign _T_4983 = _T_4153 ? 16'h2 : _T_4982; // @[Mux.scala 31:69:@2488.4]
  assign _T_4984 = _T_4150 ? 16'h1 : _T_4983; // @[Mux.scala 31:69:@2489.4]
  assign _T_4985 = _T_4984[0]; // @[OneHot.scala 66:30:@2490.4]
  assign _T_4986 = _T_4984[1]; // @[OneHot.scala 66:30:@2491.4]
  assign _T_4987 = _T_4984[2]; // @[OneHot.scala 66:30:@2492.4]
  assign _T_4988 = _T_4984[3]; // @[OneHot.scala 66:30:@2493.4]
  assign _T_4989 = _T_4984[4]; // @[OneHot.scala 66:30:@2494.4]
  assign _T_4990 = _T_4984[5]; // @[OneHot.scala 66:30:@2495.4]
  assign _T_4991 = _T_4984[6]; // @[OneHot.scala 66:30:@2496.4]
  assign _T_4992 = _T_4984[7]; // @[OneHot.scala 66:30:@2497.4]
  assign _T_4993 = _T_4984[8]; // @[OneHot.scala 66:30:@2498.4]
  assign _T_4994 = _T_4984[9]; // @[OneHot.scala 66:30:@2499.4]
  assign _T_4995 = _T_4984[10]; // @[OneHot.scala 66:30:@2500.4]
  assign _T_4996 = _T_4984[11]; // @[OneHot.scala 66:30:@2501.4]
  assign _T_4997 = _T_4984[12]; // @[OneHot.scala 66:30:@2502.4]
  assign _T_4998 = _T_4984[13]; // @[OneHot.scala 66:30:@2503.4]
  assign _T_4999 = _T_4984[14]; // @[OneHot.scala 66:30:@2504.4]
  assign _T_5000 = _T_4984[15]; // @[OneHot.scala 66:30:@2505.4]
  assign _T_5041 = _T_4150 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2523.4]
  assign _T_5042 = _T_4147 ? 16'h4000 : _T_5041; // @[Mux.scala 31:69:@2524.4]
  assign _T_5043 = _T_4144 ? 16'h2000 : _T_5042; // @[Mux.scala 31:69:@2525.4]
  assign _T_5044 = _T_4141 ? 16'h1000 : _T_5043; // @[Mux.scala 31:69:@2526.4]
  assign _T_5045 = _T_4138 ? 16'h800 : _T_5044; // @[Mux.scala 31:69:@2527.4]
  assign _T_5046 = _T_4135 ? 16'h400 : _T_5045; // @[Mux.scala 31:69:@2528.4]
  assign _T_5047 = _T_4132 ? 16'h200 : _T_5046; // @[Mux.scala 31:69:@2529.4]
  assign _T_5048 = _T_4129 ? 16'h100 : _T_5047; // @[Mux.scala 31:69:@2530.4]
  assign _T_5049 = _T_4126 ? 16'h80 : _T_5048; // @[Mux.scala 31:69:@2531.4]
  assign _T_5050 = _T_4123 ? 16'h40 : _T_5049; // @[Mux.scala 31:69:@2532.4]
  assign _T_5051 = _T_4168 ? 16'h20 : _T_5050; // @[Mux.scala 31:69:@2533.4]
  assign _T_5052 = _T_4165 ? 16'h10 : _T_5051; // @[Mux.scala 31:69:@2534.4]
  assign _T_5053 = _T_4162 ? 16'h8 : _T_5052; // @[Mux.scala 31:69:@2535.4]
  assign _T_5054 = _T_4159 ? 16'h4 : _T_5053; // @[Mux.scala 31:69:@2536.4]
  assign _T_5055 = _T_4156 ? 16'h2 : _T_5054; // @[Mux.scala 31:69:@2537.4]
  assign _T_5056 = _T_4153 ? 16'h1 : _T_5055; // @[Mux.scala 31:69:@2538.4]
  assign _T_5057 = _T_5056[0]; // @[OneHot.scala 66:30:@2539.4]
  assign _T_5058 = _T_5056[1]; // @[OneHot.scala 66:30:@2540.4]
  assign _T_5059 = _T_5056[2]; // @[OneHot.scala 66:30:@2541.4]
  assign _T_5060 = _T_5056[3]; // @[OneHot.scala 66:30:@2542.4]
  assign _T_5061 = _T_5056[4]; // @[OneHot.scala 66:30:@2543.4]
  assign _T_5062 = _T_5056[5]; // @[OneHot.scala 66:30:@2544.4]
  assign _T_5063 = _T_5056[6]; // @[OneHot.scala 66:30:@2545.4]
  assign _T_5064 = _T_5056[7]; // @[OneHot.scala 66:30:@2546.4]
  assign _T_5065 = _T_5056[8]; // @[OneHot.scala 66:30:@2547.4]
  assign _T_5066 = _T_5056[9]; // @[OneHot.scala 66:30:@2548.4]
  assign _T_5067 = _T_5056[10]; // @[OneHot.scala 66:30:@2549.4]
  assign _T_5068 = _T_5056[11]; // @[OneHot.scala 66:30:@2550.4]
  assign _T_5069 = _T_5056[12]; // @[OneHot.scala 66:30:@2551.4]
  assign _T_5070 = _T_5056[13]; // @[OneHot.scala 66:30:@2552.4]
  assign _T_5071 = _T_5056[14]; // @[OneHot.scala 66:30:@2553.4]
  assign _T_5072 = _T_5056[15]; // @[OneHot.scala 66:30:@2554.4]
  assign _T_5113 = _T_4153 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2572.4]
  assign _T_5114 = _T_4150 ? 16'h4000 : _T_5113; // @[Mux.scala 31:69:@2573.4]
  assign _T_5115 = _T_4147 ? 16'h2000 : _T_5114; // @[Mux.scala 31:69:@2574.4]
  assign _T_5116 = _T_4144 ? 16'h1000 : _T_5115; // @[Mux.scala 31:69:@2575.4]
  assign _T_5117 = _T_4141 ? 16'h800 : _T_5116; // @[Mux.scala 31:69:@2576.4]
  assign _T_5118 = _T_4138 ? 16'h400 : _T_5117; // @[Mux.scala 31:69:@2577.4]
  assign _T_5119 = _T_4135 ? 16'h200 : _T_5118; // @[Mux.scala 31:69:@2578.4]
  assign _T_5120 = _T_4132 ? 16'h100 : _T_5119; // @[Mux.scala 31:69:@2579.4]
  assign _T_5121 = _T_4129 ? 16'h80 : _T_5120; // @[Mux.scala 31:69:@2580.4]
  assign _T_5122 = _T_4126 ? 16'h40 : _T_5121; // @[Mux.scala 31:69:@2581.4]
  assign _T_5123 = _T_4123 ? 16'h20 : _T_5122; // @[Mux.scala 31:69:@2582.4]
  assign _T_5124 = _T_4168 ? 16'h10 : _T_5123; // @[Mux.scala 31:69:@2583.4]
  assign _T_5125 = _T_4165 ? 16'h8 : _T_5124; // @[Mux.scala 31:69:@2584.4]
  assign _T_5126 = _T_4162 ? 16'h4 : _T_5125; // @[Mux.scala 31:69:@2585.4]
  assign _T_5127 = _T_4159 ? 16'h2 : _T_5126; // @[Mux.scala 31:69:@2586.4]
  assign _T_5128 = _T_4156 ? 16'h1 : _T_5127; // @[Mux.scala 31:69:@2587.4]
  assign _T_5129 = _T_5128[0]; // @[OneHot.scala 66:30:@2588.4]
  assign _T_5130 = _T_5128[1]; // @[OneHot.scala 66:30:@2589.4]
  assign _T_5131 = _T_5128[2]; // @[OneHot.scala 66:30:@2590.4]
  assign _T_5132 = _T_5128[3]; // @[OneHot.scala 66:30:@2591.4]
  assign _T_5133 = _T_5128[4]; // @[OneHot.scala 66:30:@2592.4]
  assign _T_5134 = _T_5128[5]; // @[OneHot.scala 66:30:@2593.4]
  assign _T_5135 = _T_5128[6]; // @[OneHot.scala 66:30:@2594.4]
  assign _T_5136 = _T_5128[7]; // @[OneHot.scala 66:30:@2595.4]
  assign _T_5137 = _T_5128[8]; // @[OneHot.scala 66:30:@2596.4]
  assign _T_5138 = _T_5128[9]; // @[OneHot.scala 66:30:@2597.4]
  assign _T_5139 = _T_5128[10]; // @[OneHot.scala 66:30:@2598.4]
  assign _T_5140 = _T_5128[11]; // @[OneHot.scala 66:30:@2599.4]
  assign _T_5141 = _T_5128[12]; // @[OneHot.scala 66:30:@2600.4]
  assign _T_5142 = _T_5128[13]; // @[OneHot.scala 66:30:@2601.4]
  assign _T_5143 = _T_5128[14]; // @[OneHot.scala 66:30:@2602.4]
  assign _T_5144 = _T_5128[15]; // @[OneHot.scala 66:30:@2603.4]
  assign _T_5185 = _T_4156 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2621.4]
  assign _T_5186 = _T_4153 ? 16'h4000 : _T_5185; // @[Mux.scala 31:69:@2622.4]
  assign _T_5187 = _T_4150 ? 16'h2000 : _T_5186; // @[Mux.scala 31:69:@2623.4]
  assign _T_5188 = _T_4147 ? 16'h1000 : _T_5187; // @[Mux.scala 31:69:@2624.4]
  assign _T_5189 = _T_4144 ? 16'h800 : _T_5188; // @[Mux.scala 31:69:@2625.4]
  assign _T_5190 = _T_4141 ? 16'h400 : _T_5189; // @[Mux.scala 31:69:@2626.4]
  assign _T_5191 = _T_4138 ? 16'h200 : _T_5190; // @[Mux.scala 31:69:@2627.4]
  assign _T_5192 = _T_4135 ? 16'h100 : _T_5191; // @[Mux.scala 31:69:@2628.4]
  assign _T_5193 = _T_4132 ? 16'h80 : _T_5192; // @[Mux.scala 31:69:@2629.4]
  assign _T_5194 = _T_4129 ? 16'h40 : _T_5193; // @[Mux.scala 31:69:@2630.4]
  assign _T_5195 = _T_4126 ? 16'h20 : _T_5194; // @[Mux.scala 31:69:@2631.4]
  assign _T_5196 = _T_4123 ? 16'h10 : _T_5195; // @[Mux.scala 31:69:@2632.4]
  assign _T_5197 = _T_4168 ? 16'h8 : _T_5196; // @[Mux.scala 31:69:@2633.4]
  assign _T_5198 = _T_4165 ? 16'h4 : _T_5197; // @[Mux.scala 31:69:@2634.4]
  assign _T_5199 = _T_4162 ? 16'h2 : _T_5198; // @[Mux.scala 31:69:@2635.4]
  assign _T_5200 = _T_4159 ? 16'h1 : _T_5199; // @[Mux.scala 31:69:@2636.4]
  assign _T_5201 = _T_5200[0]; // @[OneHot.scala 66:30:@2637.4]
  assign _T_5202 = _T_5200[1]; // @[OneHot.scala 66:30:@2638.4]
  assign _T_5203 = _T_5200[2]; // @[OneHot.scala 66:30:@2639.4]
  assign _T_5204 = _T_5200[3]; // @[OneHot.scala 66:30:@2640.4]
  assign _T_5205 = _T_5200[4]; // @[OneHot.scala 66:30:@2641.4]
  assign _T_5206 = _T_5200[5]; // @[OneHot.scala 66:30:@2642.4]
  assign _T_5207 = _T_5200[6]; // @[OneHot.scala 66:30:@2643.4]
  assign _T_5208 = _T_5200[7]; // @[OneHot.scala 66:30:@2644.4]
  assign _T_5209 = _T_5200[8]; // @[OneHot.scala 66:30:@2645.4]
  assign _T_5210 = _T_5200[9]; // @[OneHot.scala 66:30:@2646.4]
  assign _T_5211 = _T_5200[10]; // @[OneHot.scala 66:30:@2647.4]
  assign _T_5212 = _T_5200[11]; // @[OneHot.scala 66:30:@2648.4]
  assign _T_5213 = _T_5200[12]; // @[OneHot.scala 66:30:@2649.4]
  assign _T_5214 = _T_5200[13]; // @[OneHot.scala 66:30:@2650.4]
  assign _T_5215 = _T_5200[14]; // @[OneHot.scala 66:30:@2651.4]
  assign _T_5216 = _T_5200[15]; // @[OneHot.scala 66:30:@2652.4]
  assign _T_5257 = _T_4159 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2670.4]
  assign _T_5258 = _T_4156 ? 16'h4000 : _T_5257; // @[Mux.scala 31:69:@2671.4]
  assign _T_5259 = _T_4153 ? 16'h2000 : _T_5258; // @[Mux.scala 31:69:@2672.4]
  assign _T_5260 = _T_4150 ? 16'h1000 : _T_5259; // @[Mux.scala 31:69:@2673.4]
  assign _T_5261 = _T_4147 ? 16'h800 : _T_5260; // @[Mux.scala 31:69:@2674.4]
  assign _T_5262 = _T_4144 ? 16'h400 : _T_5261; // @[Mux.scala 31:69:@2675.4]
  assign _T_5263 = _T_4141 ? 16'h200 : _T_5262; // @[Mux.scala 31:69:@2676.4]
  assign _T_5264 = _T_4138 ? 16'h100 : _T_5263; // @[Mux.scala 31:69:@2677.4]
  assign _T_5265 = _T_4135 ? 16'h80 : _T_5264; // @[Mux.scala 31:69:@2678.4]
  assign _T_5266 = _T_4132 ? 16'h40 : _T_5265; // @[Mux.scala 31:69:@2679.4]
  assign _T_5267 = _T_4129 ? 16'h20 : _T_5266; // @[Mux.scala 31:69:@2680.4]
  assign _T_5268 = _T_4126 ? 16'h10 : _T_5267; // @[Mux.scala 31:69:@2681.4]
  assign _T_5269 = _T_4123 ? 16'h8 : _T_5268; // @[Mux.scala 31:69:@2682.4]
  assign _T_5270 = _T_4168 ? 16'h4 : _T_5269; // @[Mux.scala 31:69:@2683.4]
  assign _T_5271 = _T_4165 ? 16'h2 : _T_5270; // @[Mux.scala 31:69:@2684.4]
  assign _T_5272 = _T_4162 ? 16'h1 : _T_5271; // @[Mux.scala 31:69:@2685.4]
  assign _T_5273 = _T_5272[0]; // @[OneHot.scala 66:30:@2686.4]
  assign _T_5274 = _T_5272[1]; // @[OneHot.scala 66:30:@2687.4]
  assign _T_5275 = _T_5272[2]; // @[OneHot.scala 66:30:@2688.4]
  assign _T_5276 = _T_5272[3]; // @[OneHot.scala 66:30:@2689.4]
  assign _T_5277 = _T_5272[4]; // @[OneHot.scala 66:30:@2690.4]
  assign _T_5278 = _T_5272[5]; // @[OneHot.scala 66:30:@2691.4]
  assign _T_5279 = _T_5272[6]; // @[OneHot.scala 66:30:@2692.4]
  assign _T_5280 = _T_5272[7]; // @[OneHot.scala 66:30:@2693.4]
  assign _T_5281 = _T_5272[8]; // @[OneHot.scala 66:30:@2694.4]
  assign _T_5282 = _T_5272[9]; // @[OneHot.scala 66:30:@2695.4]
  assign _T_5283 = _T_5272[10]; // @[OneHot.scala 66:30:@2696.4]
  assign _T_5284 = _T_5272[11]; // @[OneHot.scala 66:30:@2697.4]
  assign _T_5285 = _T_5272[12]; // @[OneHot.scala 66:30:@2698.4]
  assign _T_5286 = _T_5272[13]; // @[OneHot.scala 66:30:@2699.4]
  assign _T_5287 = _T_5272[14]; // @[OneHot.scala 66:30:@2700.4]
  assign _T_5288 = _T_5272[15]; // @[OneHot.scala 66:30:@2701.4]
  assign _T_5329 = _T_4162 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2719.4]
  assign _T_5330 = _T_4159 ? 16'h4000 : _T_5329; // @[Mux.scala 31:69:@2720.4]
  assign _T_5331 = _T_4156 ? 16'h2000 : _T_5330; // @[Mux.scala 31:69:@2721.4]
  assign _T_5332 = _T_4153 ? 16'h1000 : _T_5331; // @[Mux.scala 31:69:@2722.4]
  assign _T_5333 = _T_4150 ? 16'h800 : _T_5332; // @[Mux.scala 31:69:@2723.4]
  assign _T_5334 = _T_4147 ? 16'h400 : _T_5333; // @[Mux.scala 31:69:@2724.4]
  assign _T_5335 = _T_4144 ? 16'h200 : _T_5334; // @[Mux.scala 31:69:@2725.4]
  assign _T_5336 = _T_4141 ? 16'h100 : _T_5335; // @[Mux.scala 31:69:@2726.4]
  assign _T_5337 = _T_4138 ? 16'h80 : _T_5336; // @[Mux.scala 31:69:@2727.4]
  assign _T_5338 = _T_4135 ? 16'h40 : _T_5337; // @[Mux.scala 31:69:@2728.4]
  assign _T_5339 = _T_4132 ? 16'h20 : _T_5338; // @[Mux.scala 31:69:@2729.4]
  assign _T_5340 = _T_4129 ? 16'h10 : _T_5339; // @[Mux.scala 31:69:@2730.4]
  assign _T_5341 = _T_4126 ? 16'h8 : _T_5340; // @[Mux.scala 31:69:@2731.4]
  assign _T_5342 = _T_4123 ? 16'h4 : _T_5341; // @[Mux.scala 31:69:@2732.4]
  assign _T_5343 = _T_4168 ? 16'h2 : _T_5342; // @[Mux.scala 31:69:@2733.4]
  assign _T_5344 = _T_4165 ? 16'h1 : _T_5343; // @[Mux.scala 31:69:@2734.4]
  assign _T_5345 = _T_5344[0]; // @[OneHot.scala 66:30:@2735.4]
  assign _T_5346 = _T_5344[1]; // @[OneHot.scala 66:30:@2736.4]
  assign _T_5347 = _T_5344[2]; // @[OneHot.scala 66:30:@2737.4]
  assign _T_5348 = _T_5344[3]; // @[OneHot.scala 66:30:@2738.4]
  assign _T_5349 = _T_5344[4]; // @[OneHot.scala 66:30:@2739.4]
  assign _T_5350 = _T_5344[5]; // @[OneHot.scala 66:30:@2740.4]
  assign _T_5351 = _T_5344[6]; // @[OneHot.scala 66:30:@2741.4]
  assign _T_5352 = _T_5344[7]; // @[OneHot.scala 66:30:@2742.4]
  assign _T_5353 = _T_5344[8]; // @[OneHot.scala 66:30:@2743.4]
  assign _T_5354 = _T_5344[9]; // @[OneHot.scala 66:30:@2744.4]
  assign _T_5355 = _T_5344[10]; // @[OneHot.scala 66:30:@2745.4]
  assign _T_5356 = _T_5344[11]; // @[OneHot.scala 66:30:@2746.4]
  assign _T_5357 = _T_5344[12]; // @[OneHot.scala 66:30:@2747.4]
  assign _T_5358 = _T_5344[13]; // @[OneHot.scala 66:30:@2748.4]
  assign _T_5359 = _T_5344[14]; // @[OneHot.scala 66:30:@2749.4]
  assign _T_5360 = _T_5344[15]; // @[OneHot.scala 66:30:@2750.4]
  assign _T_5401 = _T_4165 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2768.4]
  assign _T_5402 = _T_4162 ? 16'h4000 : _T_5401; // @[Mux.scala 31:69:@2769.4]
  assign _T_5403 = _T_4159 ? 16'h2000 : _T_5402; // @[Mux.scala 31:69:@2770.4]
  assign _T_5404 = _T_4156 ? 16'h1000 : _T_5403; // @[Mux.scala 31:69:@2771.4]
  assign _T_5405 = _T_4153 ? 16'h800 : _T_5404; // @[Mux.scala 31:69:@2772.4]
  assign _T_5406 = _T_4150 ? 16'h400 : _T_5405; // @[Mux.scala 31:69:@2773.4]
  assign _T_5407 = _T_4147 ? 16'h200 : _T_5406; // @[Mux.scala 31:69:@2774.4]
  assign _T_5408 = _T_4144 ? 16'h100 : _T_5407; // @[Mux.scala 31:69:@2775.4]
  assign _T_5409 = _T_4141 ? 16'h80 : _T_5408; // @[Mux.scala 31:69:@2776.4]
  assign _T_5410 = _T_4138 ? 16'h40 : _T_5409; // @[Mux.scala 31:69:@2777.4]
  assign _T_5411 = _T_4135 ? 16'h20 : _T_5410; // @[Mux.scala 31:69:@2778.4]
  assign _T_5412 = _T_4132 ? 16'h10 : _T_5411; // @[Mux.scala 31:69:@2779.4]
  assign _T_5413 = _T_4129 ? 16'h8 : _T_5412; // @[Mux.scala 31:69:@2780.4]
  assign _T_5414 = _T_4126 ? 16'h4 : _T_5413; // @[Mux.scala 31:69:@2781.4]
  assign _T_5415 = _T_4123 ? 16'h2 : _T_5414; // @[Mux.scala 31:69:@2782.4]
  assign _T_5416 = _T_4168 ? 16'h1 : _T_5415; // @[Mux.scala 31:69:@2783.4]
  assign _T_5417 = _T_5416[0]; // @[OneHot.scala 66:30:@2784.4]
  assign _T_5418 = _T_5416[1]; // @[OneHot.scala 66:30:@2785.4]
  assign _T_5419 = _T_5416[2]; // @[OneHot.scala 66:30:@2786.4]
  assign _T_5420 = _T_5416[3]; // @[OneHot.scala 66:30:@2787.4]
  assign _T_5421 = _T_5416[4]; // @[OneHot.scala 66:30:@2788.4]
  assign _T_5422 = _T_5416[5]; // @[OneHot.scala 66:30:@2789.4]
  assign _T_5423 = _T_5416[6]; // @[OneHot.scala 66:30:@2790.4]
  assign _T_5424 = _T_5416[7]; // @[OneHot.scala 66:30:@2791.4]
  assign _T_5425 = _T_5416[8]; // @[OneHot.scala 66:30:@2792.4]
  assign _T_5426 = _T_5416[9]; // @[OneHot.scala 66:30:@2793.4]
  assign _T_5427 = _T_5416[10]; // @[OneHot.scala 66:30:@2794.4]
  assign _T_5428 = _T_5416[11]; // @[OneHot.scala 66:30:@2795.4]
  assign _T_5429 = _T_5416[12]; // @[OneHot.scala 66:30:@2796.4]
  assign _T_5430 = _T_5416[13]; // @[OneHot.scala 66:30:@2797.4]
  assign _T_5431 = _T_5416[14]; // @[OneHot.scala 66:30:@2798.4]
  assign _T_5432 = _T_5416[15]; // @[OneHot.scala 66:30:@2799.4]
  assign _T_5497 = {_T_4344,_T_4343,_T_4342,_T_4341,_T_4340,_T_4339,_T_4338,_T_4337}; // @[Mux.scala 19:72:@2823.4]
  assign _T_5505 = {_T_4352,_T_4351,_T_4350,_T_4349,_T_4348,_T_4347,_T_4346,_T_4345,_T_5497}; // @[Mux.scala 19:72:@2831.4]
  assign _T_5507 = _T_4265 ? _T_5505 : 16'h0; // @[Mux.scala 19:72:@2832.4]
  assign _T_5514 = {_T_4415,_T_4414,_T_4413,_T_4412,_T_4411,_T_4410,_T_4409,_T_4424}; // @[Mux.scala 19:72:@2839.4]
  assign _T_5522 = {_T_4423,_T_4422,_T_4421,_T_4420,_T_4419,_T_4418,_T_4417,_T_4416,_T_5514}; // @[Mux.scala 19:72:@2847.4]
  assign _T_5524 = _T_4266 ? _T_5522 : 16'h0; // @[Mux.scala 19:72:@2848.4]
  assign _T_5531 = {_T_4486,_T_4485,_T_4484,_T_4483,_T_4482,_T_4481,_T_4496,_T_4495}; // @[Mux.scala 19:72:@2855.4]
  assign _T_5539 = {_T_4494,_T_4493,_T_4492,_T_4491,_T_4490,_T_4489,_T_4488,_T_4487,_T_5531}; // @[Mux.scala 19:72:@2863.4]
  assign _T_5541 = _T_4267 ? _T_5539 : 16'h0; // @[Mux.scala 19:72:@2864.4]
  assign _T_5548 = {_T_4557,_T_4556,_T_4555,_T_4554,_T_4553,_T_4568,_T_4567,_T_4566}; // @[Mux.scala 19:72:@2871.4]
  assign _T_5556 = {_T_4565,_T_4564,_T_4563,_T_4562,_T_4561,_T_4560,_T_4559,_T_4558,_T_5548}; // @[Mux.scala 19:72:@2879.4]
  assign _T_5558 = _T_4268 ? _T_5556 : 16'h0; // @[Mux.scala 19:72:@2880.4]
  assign _T_5565 = {_T_4628,_T_4627,_T_4626,_T_4625,_T_4640,_T_4639,_T_4638,_T_4637}; // @[Mux.scala 19:72:@2887.4]
  assign _T_5573 = {_T_4636,_T_4635,_T_4634,_T_4633,_T_4632,_T_4631,_T_4630,_T_4629,_T_5565}; // @[Mux.scala 19:72:@2895.4]
  assign _T_5575 = _T_4269 ? _T_5573 : 16'h0; // @[Mux.scala 19:72:@2896.4]
  assign _T_5582 = {_T_4699,_T_4698,_T_4697,_T_4712,_T_4711,_T_4710,_T_4709,_T_4708}; // @[Mux.scala 19:72:@2903.4]
  assign _T_5590 = {_T_4707,_T_4706,_T_4705,_T_4704,_T_4703,_T_4702,_T_4701,_T_4700,_T_5582}; // @[Mux.scala 19:72:@2911.4]
  assign _T_5592 = _T_4270 ? _T_5590 : 16'h0; // @[Mux.scala 19:72:@2912.4]
  assign _T_5599 = {_T_4770,_T_4769,_T_4784,_T_4783,_T_4782,_T_4781,_T_4780,_T_4779}; // @[Mux.scala 19:72:@2919.4]
  assign _T_5607 = {_T_4778,_T_4777,_T_4776,_T_4775,_T_4774,_T_4773,_T_4772,_T_4771,_T_5599}; // @[Mux.scala 19:72:@2927.4]
  assign _T_5609 = _T_4271 ? _T_5607 : 16'h0; // @[Mux.scala 19:72:@2928.4]
  assign _T_5616 = {_T_4841,_T_4856,_T_4855,_T_4854,_T_4853,_T_4852,_T_4851,_T_4850}; // @[Mux.scala 19:72:@2935.4]
  assign _T_5624 = {_T_4849,_T_4848,_T_4847,_T_4846,_T_4845,_T_4844,_T_4843,_T_4842,_T_5616}; // @[Mux.scala 19:72:@2943.4]
  assign _T_5626 = _T_4272 ? _T_5624 : 16'h0; // @[Mux.scala 19:72:@2944.4]
  assign _T_5633 = {_T_4928,_T_4927,_T_4926,_T_4925,_T_4924,_T_4923,_T_4922,_T_4921}; // @[Mux.scala 19:72:@2951.4]
  assign _T_5641 = {_T_4920,_T_4919,_T_4918,_T_4917,_T_4916,_T_4915,_T_4914,_T_4913,_T_5633}; // @[Mux.scala 19:72:@2959.4]
  assign _T_5643 = _T_4273 ? _T_5641 : 16'h0; // @[Mux.scala 19:72:@2960.4]
  assign _T_5650 = {_T_4999,_T_4998,_T_4997,_T_4996,_T_4995,_T_4994,_T_4993,_T_4992}; // @[Mux.scala 19:72:@2967.4]
  assign _T_5658 = {_T_4991,_T_4990,_T_4989,_T_4988,_T_4987,_T_4986,_T_4985,_T_5000,_T_5650}; // @[Mux.scala 19:72:@2975.4]
  assign _T_5660 = _T_4274 ? _T_5658 : 16'h0; // @[Mux.scala 19:72:@2976.4]
  assign _T_5667 = {_T_5070,_T_5069,_T_5068,_T_5067,_T_5066,_T_5065,_T_5064,_T_5063}; // @[Mux.scala 19:72:@2983.4]
  assign _T_5675 = {_T_5062,_T_5061,_T_5060,_T_5059,_T_5058,_T_5057,_T_5072,_T_5071,_T_5667}; // @[Mux.scala 19:72:@2991.4]
  assign _T_5677 = _T_4275 ? _T_5675 : 16'h0; // @[Mux.scala 19:72:@2992.4]
  assign _T_5684 = {_T_5141,_T_5140,_T_5139,_T_5138,_T_5137,_T_5136,_T_5135,_T_5134}; // @[Mux.scala 19:72:@2999.4]
  assign _T_5692 = {_T_5133,_T_5132,_T_5131,_T_5130,_T_5129,_T_5144,_T_5143,_T_5142,_T_5684}; // @[Mux.scala 19:72:@3007.4]
  assign _T_5694 = _T_4276 ? _T_5692 : 16'h0; // @[Mux.scala 19:72:@3008.4]
  assign _T_5701 = {_T_5212,_T_5211,_T_5210,_T_5209,_T_5208,_T_5207,_T_5206,_T_5205}; // @[Mux.scala 19:72:@3015.4]
  assign _T_5709 = {_T_5204,_T_5203,_T_5202,_T_5201,_T_5216,_T_5215,_T_5214,_T_5213,_T_5701}; // @[Mux.scala 19:72:@3023.4]
  assign _T_5711 = _T_4277 ? _T_5709 : 16'h0; // @[Mux.scala 19:72:@3024.4]
  assign _T_5718 = {_T_5283,_T_5282,_T_5281,_T_5280,_T_5279,_T_5278,_T_5277,_T_5276}; // @[Mux.scala 19:72:@3031.4]
  assign _T_5726 = {_T_5275,_T_5274,_T_5273,_T_5288,_T_5287,_T_5286,_T_5285,_T_5284,_T_5718}; // @[Mux.scala 19:72:@3039.4]
  assign _T_5728 = _T_4278 ? _T_5726 : 16'h0; // @[Mux.scala 19:72:@3040.4]
  assign _T_5735 = {_T_5354,_T_5353,_T_5352,_T_5351,_T_5350,_T_5349,_T_5348,_T_5347}; // @[Mux.scala 19:72:@3047.4]
  assign _T_5743 = {_T_5346,_T_5345,_T_5360,_T_5359,_T_5358,_T_5357,_T_5356,_T_5355,_T_5735}; // @[Mux.scala 19:72:@3055.4]
  assign _T_5745 = _T_4279 ? _T_5743 : 16'h0; // @[Mux.scala 19:72:@3056.4]
  assign _T_5752 = {_T_5425,_T_5424,_T_5423,_T_5422,_T_5421,_T_5420,_T_5419,_T_5418}; // @[Mux.scala 19:72:@3063.4]
  assign _T_5760 = {_T_5417,_T_5432,_T_5431,_T_5430,_T_5429,_T_5428,_T_5427,_T_5426,_T_5752}; // @[Mux.scala 19:72:@3071.4]
  assign _T_5762 = _T_4280 ? _T_5760 : 16'h0; // @[Mux.scala 19:72:@3072.4]
  assign _T_5763 = _T_5507 | _T_5524; // @[Mux.scala 19:72:@3073.4]
  assign _T_5764 = _T_5763 | _T_5541; // @[Mux.scala 19:72:@3074.4]
  assign _T_5765 = _T_5764 | _T_5558; // @[Mux.scala 19:72:@3075.4]
  assign _T_5766 = _T_5765 | _T_5575; // @[Mux.scala 19:72:@3076.4]
  assign _T_5767 = _T_5766 | _T_5592; // @[Mux.scala 19:72:@3077.4]
  assign _T_5768 = _T_5767 | _T_5609; // @[Mux.scala 19:72:@3078.4]
  assign _T_5769 = _T_5768 | _T_5626; // @[Mux.scala 19:72:@3079.4]
  assign _T_5770 = _T_5769 | _T_5643; // @[Mux.scala 19:72:@3080.4]
  assign _T_5771 = _T_5770 | _T_5660; // @[Mux.scala 19:72:@3081.4]
  assign _T_5772 = _T_5771 | _T_5677; // @[Mux.scala 19:72:@3082.4]
  assign _T_5773 = _T_5772 | _T_5694; // @[Mux.scala 19:72:@3083.4]
  assign _T_5774 = _T_5773 | _T_5711; // @[Mux.scala 19:72:@3084.4]
  assign _T_5775 = _T_5774 | _T_5728; // @[Mux.scala 19:72:@3085.4]
  assign _T_5776 = _T_5775 | _T_5745; // @[Mux.scala 19:72:@3086.4]
  assign _T_5777 = _T_5776 | _T_5762; // @[Mux.scala 19:72:@3087.4]
  assign inputAddrPriorityPorts_0_0 = _T_5777[0]; // @[Mux.scala 19:72:@3091.4]
  assign inputAddrPriorityPorts_0_1 = _T_5777[1]; // @[Mux.scala 19:72:@3093.4]
  assign inputAddrPriorityPorts_0_2 = _T_5777[2]; // @[Mux.scala 19:72:@3095.4]
  assign inputAddrPriorityPorts_0_3 = _T_5777[3]; // @[Mux.scala 19:72:@3097.4]
  assign inputAddrPriorityPorts_0_4 = _T_5777[4]; // @[Mux.scala 19:72:@3099.4]
  assign inputAddrPriorityPorts_0_5 = _T_5777[5]; // @[Mux.scala 19:72:@3101.4]
  assign inputAddrPriorityPorts_0_6 = _T_5777[6]; // @[Mux.scala 19:72:@3103.4]
  assign inputAddrPriorityPorts_0_7 = _T_5777[7]; // @[Mux.scala 19:72:@3105.4]
  assign inputAddrPriorityPorts_0_8 = _T_5777[8]; // @[Mux.scala 19:72:@3107.4]
  assign inputAddrPriorityPorts_0_9 = _T_5777[9]; // @[Mux.scala 19:72:@3109.4]
  assign inputAddrPriorityPorts_0_10 = _T_5777[10]; // @[Mux.scala 19:72:@3111.4]
  assign inputAddrPriorityPorts_0_11 = _T_5777[11]; // @[Mux.scala 19:72:@3113.4]
  assign inputAddrPriorityPorts_0_12 = _T_5777[12]; // @[Mux.scala 19:72:@3115.4]
  assign inputAddrPriorityPorts_0_13 = _T_5777[13]; // @[Mux.scala 19:72:@3117.4]
  assign inputAddrPriorityPorts_0_14 = _T_5777[14]; // @[Mux.scala 19:72:@3119.4]
  assign inputAddrPriorityPorts_0_15 = _T_5777[15]; // @[Mux.scala 19:72:@3121.4]
  assign _T_5979 = _T_4238 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3175.4]
  assign _T_5980 = _T_4235 ? 16'h4000 : _T_5979; // @[Mux.scala 31:69:@3176.4]
  assign _T_5981 = _T_4232 ? 16'h2000 : _T_5980; // @[Mux.scala 31:69:@3177.4]
  assign _T_5982 = _T_4229 ? 16'h1000 : _T_5981; // @[Mux.scala 31:69:@3178.4]
  assign _T_5983 = _T_4226 ? 16'h800 : _T_5982; // @[Mux.scala 31:69:@3179.4]
  assign _T_5984 = _T_4223 ? 16'h400 : _T_5983; // @[Mux.scala 31:69:@3180.4]
  assign _T_5985 = _T_4220 ? 16'h200 : _T_5984; // @[Mux.scala 31:69:@3181.4]
  assign _T_5986 = _T_4217 ? 16'h100 : _T_5985; // @[Mux.scala 31:69:@3182.4]
  assign _T_5987 = _T_4214 ? 16'h80 : _T_5986; // @[Mux.scala 31:69:@3183.4]
  assign _T_5988 = _T_4211 ? 16'h40 : _T_5987; // @[Mux.scala 31:69:@3184.4]
  assign _T_5989 = _T_4208 ? 16'h20 : _T_5988; // @[Mux.scala 31:69:@3185.4]
  assign _T_5990 = _T_4205 ? 16'h10 : _T_5989; // @[Mux.scala 31:69:@3186.4]
  assign _T_5991 = _T_4202 ? 16'h8 : _T_5990; // @[Mux.scala 31:69:@3187.4]
  assign _T_5992 = _T_4199 ? 16'h4 : _T_5991; // @[Mux.scala 31:69:@3188.4]
  assign _T_5993 = _T_4196 ? 16'h2 : _T_5992; // @[Mux.scala 31:69:@3189.4]
  assign _T_5994 = _T_4193 ? 16'h1 : _T_5993; // @[Mux.scala 31:69:@3190.4]
  assign _T_5995 = _T_5994[0]; // @[OneHot.scala 66:30:@3191.4]
  assign _T_5996 = _T_5994[1]; // @[OneHot.scala 66:30:@3192.4]
  assign _T_5997 = _T_5994[2]; // @[OneHot.scala 66:30:@3193.4]
  assign _T_5998 = _T_5994[3]; // @[OneHot.scala 66:30:@3194.4]
  assign _T_5999 = _T_5994[4]; // @[OneHot.scala 66:30:@3195.4]
  assign _T_6000 = _T_5994[5]; // @[OneHot.scala 66:30:@3196.4]
  assign _T_6001 = _T_5994[6]; // @[OneHot.scala 66:30:@3197.4]
  assign _T_6002 = _T_5994[7]; // @[OneHot.scala 66:30:@3198.4]
  assign _T_6003 = _T_5994[8]; // @[OneHot.scala 66:30:@3199.4]
  assign _T_6004 = _T_5994[9]; // @[OneHot.scala 66:30:@3200.4]
  assign _T_6005 = _T_5994[10]; // @[OneHot.scala 66:30:@3201.4]
  assign _T_6006 = _T_5994[11]; // @[OneHot.scala 66:30:@3202.4]
  assign _T_6007 = _T_5994[12]; // @[OneHot.scala 66:30:@3203.4]
  assign _T_6008 = _T_5994[13]; // @[OneHot.scala 66:30:@3204.4]
  assign _T_6009 = _T_5994[14]; // @[OneHot.scala 66:30:@3205.4]
  assign _T_6010 = _T_5994[15]; // @[OneHot.scala 66:30:@3206.4]
  assign _T_6051 = _T_4193 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3224.4]
  assign _T_6052 = _T_4238 ? 16'h4000 : _T_6051; // @[Mux.scala 31:69:@3225.4]
  assign _T_6053 = _T_4235 ? 16'h2000 : _T_6052; // @[Mux.scala 31:69:@3226.4]
  assign _T_6054 = _T_4232 ? 16'h1000 : _T_6053; // @[Mux.scala 31:69:@3227.4]
  assign _T_6055 = _T_4229 ? 16'h800 : _T_6054; // @[Mux.scala 31:69:@3228.4]
  assign _T_6056 = _T_4226 ? 16'h400 : _T_6055; // @[Mux.scala 31:69:@3229.4]
  assign _T_6057 = _T_4223 ? 16'h200 : _T_6056; // @[Mux.scala 31:69:@3230.4]
  assign _T_6058 = _T_4220 ? 16'h100 : _T_6057; // @[Mux.scala 31:69:@3231.4]
  assign _T_6059 = _T_4217 ? 16'h80 : _T_6058; // @[Mux.scala 31:69:@3232.4]
  assign _T_6060 = _T_4214 ? 16'h40 : _T_6059; // @[Mux.scala 31:69:@3233.4]
  assign _T_6061 = _T_4211 ? 16'h20 : _T_6060; // @[Mux.scala 31:69:@3234.4]
  assign _T_6062 = _T_4208 ? 16'h10 : _T_6061; // @[Mux.scala 31:69:@3235.4]
  assign _T_6063 = _T_4205 ? 16'h8 : _T_6062; // @[Mux.scala 31:69:@3236.4]
  assign _T_6064 = _T_4202 ? 16'h4 : _T_6063; // @[Mux.scala 31:69:@3237.4]
  assign _T_6065 = _T_4199 ? 16'h2 : _T_6064; // @[Mux.scala 31:69:@3238.4]
  assign _T_6066 = _T_4196 ? 16'h1 : _T_6065; // @[Mux.scala 31:69:@3239.4]
  assign _T_6067 = _T_6066[0]; // @[OneHot.scala 66:30:@3240.4]
  assign _T_6068 = _T_6066[1]; // @[OneHot.scala 66:30:@3241.4]
  assign _T_6069 = _T_6066[2]; // @[OneHot.scala 66:30:@3242.4]
  assign _T_6070 = _T_6066[3]; // @[OneHot.scala 66:30:@3243.4]
  assign _T_6071 = _T_6066[4]; // @[OneHot.scala 66:30:@3244.4]
  assign _T_6072 = _T_6066[5]; // @[OneHot.scala 66:30:@3245.4]
  assign _T_6073 = _T_6066[6]; // @[OneHot.scala 66:30:@3246.4]
  assign _T_6074 = _T_6066[7]; // @[OneHot.scala 66:30:@3247.4]
  assign _T_6075 = _T_6066[8]; // @[OneHot.scala 66:30:@3248.4]
  assign _T_6076 = _T_6066[9]; // @[OneHot.scala 66:30:@3249.4]
  assign _T_6077 = _T_6066[10]; // @[OneHot.scala 66:30:@3250.4]
  assign _T_6078 = _T_6066[11]; // @[OneHot.scala 66:30:@3251.4]
  assign _T_6079 = _T_6066[12]; // @[OneHot.scala 66:30:@3252.4]
  assign _T_6080 = _T_6066[13]; // @[OneHot.scala 66:30:@3253.4]
  assign _T_6081 = _T_6066[14]; // @[OneHot.scala 66:30:@3254.4]
  assign _T_6082 = _T_6066[15]; // @[OneHot.scala 66:30:@3255.4]
  assign _T_6123 = _T_4196 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3273.4]
  assign _T_6124 = _T_4193 ? 16'h4000 : _T_6123; // @[Mux.scala 31:69:@3274.4]
  assign _T_6125 = _T_4238 ? 16'h2000 : _T_6124; // @[Mux.scala 31:69:@3275.4]
  assign _T_6126 = _T_4235 ? 16'h1000 : _T_6125; // @[Mux.scala 31:69:@3276.4]
  assign _T_6127 = _T_4232 ? 16'h800 : _T_6126; // @[Mux.scala 31:69:@3277.4]
  assign _T_6128 = _T_4229 ? 16'h400 : _T_6127; // @[Mux.scala 31:69:@3278.4]
  assign _T_6129 = _T_4226 ? 16'h200 : _T_6128; // @[Mux.scala 31:69:@3279.4]
  assign _T_6130 = _T_4223 ? 16'h100 : _T_6129; // @[Mux.scala 31:69:@3280.4]
  assign _T_6131 = _T_4220 ? 16'h80 : _T_6130; // @[Mux.scala 31:69:@3281.4]
  assign _T_6132 = _T_4217 ? 16'h40 : _T_6131; // @[Mux.scala 31:69:@3282.4]
  assign _T_6133 = _T_4214 ? 16'h20 : _T_6132; // @[Mux.scala 31:69:@3283.4]
  assign _T_6134 = _T_4211 ? 16'h10 : _T_6133; // @[Mux.scala 31:69:@3284.4]
  assign _T_6135 = _T_4208 ? 16'h8 : _T_6134; // @[Mux.scala 31:69:@3285.4]
  assign _T_6136 = _T_4205 ? 16'h4 : _T_6135; // @[Mux.scala 31:69:@3286.4]
  assign _T_6137 = _T_4202 ? 16'h2 : _T_6136; // @[Mux.scala 31:69:@3287.4]
  assign _T_6138 = _T_4199 ? 16'h1 : _T_6137; // @[Mux.scala 31:69:@3288.4]
  assign _T_6139 = _T_6138[0]; // @[OneHot.scala 66:30:@3289.4]
  assign _T_6140 = _T_6138[1]; // @[OneHot.scala 66:30:@3290.4]
  assign _T_6141 = _T_6138[2]; // @[OneHot.scala 66:30:@3291.4]
  assign _T_6142 = _T_6138[3]; // @[OneHot.scala 66:30:@3292.4]
  assign _T_6143 = _T_6138[4]; // @[OneHot.scala 66:30:@3293.4]
  assign _T_6144 = _T_6138[5]; // @[OneHot.scala 66:30:@3294.4]
  assign _T_6145 = _T_6138[6]; // @[OneHot.scala 66:30:@3295.4]
  assign _T_6146 = _T_6138[7]; // @[OneHot.scala 66:30:@3296.4]
  assign _T_6147 = _T_6138[8]; // @[OneHot.scala 66:30:@3297.4]
  assign _T_6148 = _T_6138[9]; // @[OneHot.scala 66:30:@3298.4]
  assign _T_6149 = _T_6138[10]; // @[OneHot.scala 66:30:@3299.4]
  assign _T_6150 = _T_6138[11]; // @[OneHot.scala 66:30:@3300.4]
  assign _T_6151 = _T_6138[12]; // @[OneHot.scala 66:30:@3301.4]
  assign _T_6152 = _T_6138[13]; // @[OneHot.scala 66:30:@3302.4]
  assign _T_6153 = _T_6138[14]; // @[OneHot.scala 66:30:@3303.4]
  assign _T_6154 = _T_6138[15]; // @[OneHot.scala 66:30:@3304.4]
  assign _T_6195 = _T_4199 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3322.4]
  assign _T_6196 = _T_4196 ? 16'h4000 : _T_6195; // @[Mux.scala 31:69:@3323.4]
  assign _T_6197 = _T_4193 ? 16'h2000 : _T_6196; // @[Mux.scala 31:69:@3324.4]
  assign _T_6198 = _T_4238 ? 16'h1000 : _T_6197; // @[Mux.scala 31:69:@3325.4]
  assign _T_6199 = _T_4235 ? 16'h800 : _T_6198; // @[Mux.scala 31:69:@3326.4]
  assign _T_6200 = _T_4232 ? 16'h400 : _T_6199; // @[Mux.scala 31:69:@3327.4]
  assign _T_6201 = _T_4229 ? 16'h200 : _T_6200; // @[Mux.scala 31:69:@3328.4]
  assign _T_6202 = _T_4226 ? 16'h100 : _T_6201; // @[Mux.scala 31:69:@3329.4]
  assign _T_6203 = _T_4223 ? 16'h80 : _T_6202; // @[Mux.scala 31:69:@3330.4]
  assign _T_6204 = _T_4220 ? 16'h40 : _T_6203; // @[Mux.scala 31:69:@3331.4]
  assign _T_6205 = _T_4217 ? 16'h20 : _T_6204; // @[Mux.scala 31:69:@3332.4]
  assign _T_6206 = _T_4214 ? 16'h10 : _T_6205; // @[Mux.scala 31:69:@3333.4]
  assign _T_6207 = _T_4211 ? 16'h8 : _T_6206; // @[Mux.scala 31:69:@3334.4]
  assign _T_6208 = _T_4208 ? 16'h4 : _T_6207; // @[Mux.scala 31:69:@3335.4]
  assign _T_6209 = _T_4205 ? 16'h2 : _T_6208; // @[Mux.scala 31:69:@3336.4]
  assign _T_6210 = _T_4202 ? 16'h1 : _T_6209; // @[Mux.scala 31:69:@3337.4]
  assign _T_6211 = _T_6210[0]; // @[OneHot.scala 66:30:@3338.4]
  assign _T_6212 = _T_6210[1]; // @[OneHot.scala 66:30:@3339.4]
  assign _T_6213 = _T_6210[2]; // @[OneHot.scala 66:30:@3340.4]
  assign _T_6214 = _T_6210[3]; // @[OneHot.scala 66:30:@3341.4]
  assign _T_6215 = _T_6210[4]; // @[OneHot.scala 66:30:@3342.4]
  assign _T_6216 = _T_6210[5]; // @[OneHot.scala 66:30:@3343.4]
  assign _T_6217 = _T_6210[6]; // @[OneHot.scala 66:30:@3344.4]
  assign _T_6218 = _T_6210[7]; // @[OneHot.scala 66:30:@3345.4]
  assign _T_6219 = _T_6210[8]; // @[OneHot.scala 66:30:@3346.4]
  assign _T_6220 = _T_6210[9]; // @[OneHot.scala 66:30:@3347.4]
  assign _T_6221 = _T_6210[10]; // @[OneHot.scala 66:30:@3348.4]
  assign _T_6222 = _T_6210[11]; // @[OneHot.scala 66:30:@3349.4]
  assign _T_6223 = _T_6210[12]; // @[OneHot.scala 66:30:@3350.4]
  assign _T_6224 = _T_6210[13]; // @[OneHot.scala 66:30:@3351.4]
  assign _T_6225 = _T_6210[14]; // @[OneHot.scala 66:30:@3352.4]
  assign _T_6226 = _T_6210[15]; // @[OneHot.scala 66:30:@3353.4]
  assign _T_6267 = _T_4202 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3371.4]
  assign _T_6268 = _T_4199 ? 16'h4000 : _T_6267; // @[Mux.scala 31:69:@3372.4]
  assign _T_6269 = _T_4196 ? 16'h2000 : _T_6268; // @[Mux.scala 31:69:@3373.4]
  assign _T_6270 = _T_4193 ? 16'h1000 : _T_6269; // @[Mux.scala 31:69:@3374.4]
  assign _T_6271 = _T_4238 ? 16'h800 : _T_6270; // @[Mux.scala 31:69:@3375.4]
  assign _T_6272 = _T_4235 ? 16'h400 : _T_6271; // @[Mux.scala 31:69:@3376.4]
  assign _T_6273 = _T_4232 ? 16'h200 : _T_6272; // @[Mux.scala 31:69:@3377.4]
  assign _T_6274 = _T_4229 ? 16'h100 : _T_6273; // @[Mux.scala 31:69:@3378.4]
  assign _T_6275 = _T_4226 ? 16'h80 : _T_6274; // @[Mux.scala 31:69:@3379.4]
  assign _T_6276 = _T_4223 ? 16'h40 : _T_6275; // @[Mux.scala 31:69:@3380.4]
  assign _T_6277 = _T_4220 ? 16'h20 : _T_6276; // @[Mux.scala 31:69:@3381.4]
  assign _T_6278 = _T_4217 ? 16'h10 : _T_6277; // @[Mux.scala 31:69:@3382.4]
  assign _T_6279 = _T_4214 ? 16'h8 : _T_6278; // @[Mux.scala 31:69:@3383.4]
  assign _T_6280 = _T_4211 ? 16'h4 : _T_6279; // @[Mux.scala 31:69:@3384.4]
  assign _T_6281 = _T_4208 ? 16'h2 : _T_6280; // @[Mux.scala 31:69:@3385.4]
  assign _T_6282 = _T_4205 ? 16'h1 : _T_6281; // @[Mux.scala 31:69:@3386.4]
  assign _T_6283 = _T_6282[0]; // @[OneHot.scala 66:30:@3387.4]
  assign _T_6284 = _T_6282[1]; // @[OneHot.scala 66:30:@3388.4]
  assign _T_6285 = _T_6282[2]; // @[OneHot.scala 66:30:@3389.4]
  assign _T_6286 = _T_6282[3]; // @[OneHot.scala 66:30:@3390.4]
  assign _T_6287 = _T_6282[4]; // @[OneHot.scala 66:30:@3391.4]
  assign _T_6288 = _T_6282[5]; // @[OneHot.scala 66:30:@3392.4]
  assign _T_6289 = _T_6282[6]; // @[OneHot.scala 66:30:@3393.4]
  assign _T_6290 = _T_6282[7]; // @[OneHot.scala 66:30:@3394.4]
  assign _T_6291 = _T_6282[8]; // @[OneHot.scala 66:30:@3395.4]
  assign _T_6292 = _T_6282[9]; // @[OneHot.scala 66:30:@3396.4]
  assign _T_6293 = _T_6282[10]; // @[OneHot.scala 66:30:@3397.4]
  assign _T_6294 = _T_6282[11]; // @[OneHot.scala 66:30:@3398.4]
  assign _T_6295 = _T_6282[12]; // @[OneHot.scala 66:30:@3399.4]
  assign _T_6296 = _T_6282[13]; // @[OneHot.scala 66:30:@3400.4]
  assign _T_6297 = _T_6282[14]; // @[OneHot.scala 66:30:@3401.4]
  assign _T_6298 = _T_6282[15]; // @[OneHot.scala 66:30:@3402.4]
  assign _T_6339 = _T_4205 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3420.4]
  assign _T_6340 = _T_4202 ? 16'h4000 : _T_6339; // @[Mux.scala 31:69:@3421.4]
  assign _T_6341 = _T_4199 ? 16'h2000 : _T_6340; // @[Mux.scala 31:69:@3422.4]
  assign _T_6342 = _T_4196 ? 16'h1000 : _T_6341; // @[Mux.scala 31:69:@3423.4]
  assign _T_6343 = _T_4193 ? 16'h800 : _T_6342; // @[Mux.scala 31:69:@3424.4]
  assign _T_6344 = _T_4238 ? 16'h400 : _T_6343; // @[Mux.scala 31:69:@3425.4]
  assign _T_6345 = _T_4235 ? 16'h200 : _T_6344; // @[Mux.scala 31:69:@3426.4]
  assign _T_6346 = _T_4232 ? 16'h100 : _T_6345; // @[Mux.scala 31:69:@3427.4]
  assign _T_6347 = _T_4229 ? 16'h80 : _T_6346; // @[Mux.scala 31:69:@3428.4]
  assign _T_6348 = _T_4226 ? 16'h40 : _T_6347; // @[Mux.scala 31:69:@3429.4]
  assign _T_6349 = _T_4223 ? 16'h20 : _T_6348; // @[Mux.scala 31:69:@3430.4]
  assign _T_6350 = _T_4220 ? 16'h10 : _T_6349; // @[Mux.scala 31:69:@3431.4]
  assign _T_6351 = _T_4217 ? 16'h8 : _T_6350; // @[Mux.scala 31:69:@3432.4]
  assign _T_6352 = _T_4214 ? 16'h4 : _T_6351; // @[Mux.scala 31:69:@3433.4]
  assign _T_6353 = _T_4211 ? 16'h2 : _T_6352; // @[Mux.scala 31:69:@3434.4]
  assign _T_6354 = _T_4208 ? 16'h1 : _T_6353; // @[Mux.scala 31:69:@3435.4]
  assign _T_6355 = _T_6354[0]; // @[OneHot.scala 66:30:@3436.4]
  assign _T_6356 = _T_6354[1]; // @[OneHot.scala 66:30:@3437.4]
  assign _T_6357 = _T_6354[2]; // @[OneHot.scala 66:30:@3438.4]
  assign _T_6358 = _T_6354[3]; // @[OneHot.scala 66:30:@3439.4]
  assign _T_6359 = _T_6354[4]; // @[OneHot.scala 66:30:@3440.4]
  assign _T_6360 = _T_6354[5]; // @[OneHot.scala 66:30:@3441.4]
  assign _T_6361 = _T_6354[6]; // @[OneHot.scala 66:30:@3442.4]
  assign _T_6362 = _T_6354[7]; // @[OneHot.scala 66:30:@3443.4]
  assign _T_6363 = _T_6354[8]; // @[OneHot.scala 66:30:@3444.4]
  assign _T_6364 = _T_6354[9]; // @[OneHot.scala 66:30:@3445.4]
  assign _T_6365 = _T_6354[10]; // @[OneHot.scala 66:30:@3446.4]
  assign _T_6366 = _T_6354[11]; // @[OneHot.scala 66:30:@3447.4]
  assign _T_6367 = _T_6354[12]; // @[OneHot.scala 66:30:@3448.4]
  assign _T_6368 = _T_6354[13]; // @[OneHot.scala 66:30:@3449.4]
  assign _T_6369 = _T_6354[14]; // @[OneHot.scala 66:30:@3450.4]
  assign _T_6370 = _T_6354[15]; // @[OneHot.scala 66:30:@3451.4]
  assign _T_6411 = _T_4208 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3469.4]
  assign _T_6412 = _T_4205 ? 16'h4000 : _T_6411; // @[Mux.scala 31:69:@3470.4]
  assign _T_6413 = _T_4202 ? 16'h2000 : _T_6412; // @[Mux.scala 31:69:@3471.4]
  assign _T_6414 = _T_4199 ? 16'h1000 : _T_6413; // @[Mux.scala 31:69:@3472.4]
  assign _T_6415 = _T_4196 ? 16'h800 : _T_6414; // @[Mux.scala 31:69:@3473.4]
  assign _T_6416 = _T_4193 ? 16'h400 : _T_6415; // @[Mux.scala 31:69:@3474.4]
  assign _T_6417 = _T_4238 ? 16'h200 : _T_6416; // @[Mux.scala 31:69:@3475.4]
  assign _T_6418 = _T_4235 ? 16'h100 : _T_6417; // @[Mux.scala 31:69:@3476.4]
  assign _T_6419 = _T_4232 ? 16'h80 : _T_6418; // @[Mux.scala 31:69:@3477.4]
  assign _T_6420 = _T_4229 ? 16'h40 : _T_6419; // @[Mux.scala 31:69:@3478.4]
  assign _T_6421 = _T_4226 ? 16'h20 : _T_6420; // @[Mux.scala 31:69:@3479.4]
  assign _T_6422 = _T_4223 ? 16'h10 : _T_6421; // @[Mux.scala 31:69:@3480.4]
  assign _T_6423 = _T_4220 ? 16'h8 : _T_6422; // @[Mux.scala 31:69:@3481.4]
  assign _T_6424 = _T_4217 ? 16'h4 : _T_6423; // @[Mux.scala 31:69:@3482.4]
  assign _T_6425 = _T_4214 ? 16'h2 : _T_6424; // @[Mux.scala 31:69:@3483.4]
  assign _T_6426 = _T_4211 ? 16'h1 : _T_6425; // @[Mux.scala 31:69:@3484.4]
  assign _T_6427 = _T_6426[0]; // @[OneHot.scala 66:30:@3485.4]
  assign _T_6428 = _T_6426[1]; // @[OneHot.scala 66:30:@3486.4]
  assign _T_6429 = _T_6426[2]; // @[OneHot.scala 66:30:@3487.4]
  assign _T_6430 = _T_6426[3]; // @[OneHot.scala 66:30:@3488.4]
  assign _T_6431 = _T_6426[4]; // @[OneHot.scala 66:30:@3489.4]
  assign _T_6432 = _T_6426[5]; // @[OneHot.scala 66:30:@3490.4]
  assign _T_6433 = _T_6426[6]; // @[OneHot.scala 66:30:@3491.4]
  assign _T_6434 = _T_6426[7]; // @[OneHot.scala 66:30:@3492.4]
  assign _T_6435 = _T_6426[8]; // @[OneHot.scala 66:30:@3493.4]
  assign _T_6436 = _T_6426[9]; // @[OneHot.scala 66:30:@3494.4]
  assign _T_6437 = _T_6426[10]; // @[OneHot.scala 66:30:@3495.4]
  assign _T_6438 = _T_6426[11]; // @[OneHot.scala 66:30:@3496.4]
  assign _T_6439 = _T_6426[12]; // @[OneHot.scala 66:30:@3497.4]
  assign _T_6440 = _T_6426[13]; // @[OneHot.scala 66:30:@3498.4]
  assign _T_6441 = _T_6426[14]; // @[OneHot.scala 66:30:@3499.4]
  assign _T_6442 = _T_6426[15]; // @[OneHot.scala 66:30:@3500.4]
  assign _T_6483 = _T_4211 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3518.4]
  assign _T_6484 = _T_4208 ? 16'h4000 : _T_6483; // @[Mux.scala 31:69:@3519.4]
  assign _T_6485 = _T_4205 ? 16'h2000 : _T_6484; // @[Mux.scala 31:69:@3520.4]
  assign _T_6486 = _T_4202 ? 16'h1000 : _T_6485; // @[Mux.scala 31:69:@3521.4]
  assign _T_6487 = _T_4199 ? 16'h800 : _T_6486; // @[Mux.scala 31:69:@3522.4]
  assign _T_6488 = _T_4196 ? 16'h400 : _T_6487; // @[Mux.scala 31:69:@3523.4]
  assign _T_6489 = _T_4193 ? 16'h200 : _T_6488; // @[Mux.scala 31:69:@3524.4]
  assign _T_6490 = _T_4238 ? 16'h100 : _T_6489; // @[Mux.scala 31:69:@3525.4]
  assign _T_6491 = _T_4235 ? 16'h80 : _T_6490; // @[Mux.scala 31:69:@3526.4]
  assign _T_6492 = _T_4232 ? 16'h40 : _T_6491; // @[Mux.scala 31:69:@3527.4]
  assign _T_6493 = _T_4229 ? 16'h20 : _T_6492; // @[Mux.scala 31:69:@3528.4]
  assign _T_6494 = _T_4226 ? 16'h10 : _T_6493; // @[Mux.scala 31:69:@3529.4]
  assign _T_6495 = _T_4223 ? 16'h8 : _T_6494; // @[Mux.scala 31:69:@3530.4]
  assign _T_6496 = _T_4220 ? 16'h4 : _T_6495; // @[Mux.scala 31:69:@3531.4]
  assign _T_6497 = _T_4217 ? 16'h2 : _T_6496; // @[Mux.scala 31:69:@3532.4]
  assign _T_6498 = _T_4214 ? 16'h1 : _T_6497; // @[Mux.scala 31:69:@3533.4]
  assign _T_6499 = _T_6498[0]; // @[OneHot.scala 66:30:@3534.4]
  assign _T_6500 = _T_6498[1]; // @[OneHot.scala 66:30:@3535.4]
  assign _T_6501 = _T_6498[2]; // @[OneHot.scala 66:30:@3536.4]
  assign _T_6502 = _T_6498[3]; // @[OneHot.scala 66:30:@3537.4]
  assign _T_6503 = _T_6498[4]; // @[OneHot.scala 66:30:@3538.4]
  assign _T_6504 = _T_6498[5]; // @[OneHot.scala 66:30:@3539.4]
  assign _T_6505 = _T_6498[6]; // @[OneHot.scala 66:30:@3540.4]
  assign _T_6506 = _T_6498[7]; // @[OneHot.scala 66:30:@3541.4]
  assign _T_6507 = _T_6498[8]; // @[OneHot.scala 66:30:@3542.4]
  assign _T_6508 = _T_6498[9]; // @[OneHot.scala 66:30:@3543.4]
  assign _T_6509 = _T_6498[10]; // @[OneHot.scala 66:30:@3544.4]
  assign _T_6510 = _T_6498[11]; // @[OneHot.scala 66:30:@3545.4]
  assign _T_6511 = _T_6498[12]; // @[OneHot.scala 66:30:@3546.4]
  assign _T_6512 = _T_6498[13]; // @[OneHot.scala 66:30:@3547.4]
  assign _T_6513 = _T_6498[14]; // @[OneHot.scala 66:30:@3548.4]
  assign _T_6514 = _T_6498[15]; // @[OneHot.scala 66:30:@3549.4]
  assign _T_6555 = _T_4214 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3567.4]
  assign _T_6556 = _T_4211 ? 16'h4000 : _T_6555; // @[Mux.scala 31:69:@3568.4]
  assign _T_6557 = _T_4208 ? 16'h2000 : _T_6556; // @[Mux.scala 31:69:@3569.4]
  assign _T_6558 = _T_4205 ? 16'h1000 : _T_6557; // @[Mux.scala 31:69:@3570.4]
  assign _T_6559 = _T_4202 ? 16'h800 : _T_6558; // @[Mux.scala 31:69:@3571.4]
  assign _T_6560 = _T_4199 ? 16'h400 : _T_6559; // @[Mux.scala 31:69:@3572.4]
  assign _T_6561 = _T_4196 ? 16'h200 : _T_6560; // @[Mux.scala 31:69:@3573.4]
  assign _T_6562 = _T_4193 ? 16'h100 : _T_6561; // @[Mux.scala 31:69:@3574.4]
  assign _T_6563 = _T_4238 ? 16'h80 : _T_6562; // @[Mux.scala 31:69:@3575.4]
  assign _T_6564 = _T_4235 ? 16'h40 : _T_6563; // @[Mux.scala 31:69:@3576.4]
  assign _T_6565 = _T_4232 ? 16'h20 : _T_6564; // @[Mux.scala 31:69:@3577.4]
  assign _T_6566 = _T_4229 ? 16'h10 : _T_6565; // @[Mux.scala 31:69:@3578.4]
  assign _T_6567 = _T_4226 ? 16'h8 : _T_6566; // @[Mux.scala 31:69:@3579.4]
  assign _T_6568 = _T_4223 ? 16'h4 : _T_6567; // @[Mux.scala 31:69:@3580.4]
  assign _T_6569 = _T_4220 ? 16'h2 : _T_6568; // @[Mux.scala 31:69:@3581.4]
  assign _T_6570 = _T_4217 ? 16'h1 : _T_6569; // @[Mux.scala 31:69:@3582.4]
  assign _T_6571 = _T_6570[0]; // @[OneHot.scala 66:30:@3583.4]
  assign _T_6572 = _T_6570[1]; // @[OneHot.scala 66:30:@3584.4]
  assign _T_6573 = _T_6570[2]; // @[OneHot.scala 66:30:@3585.4]
  assign _T_6574 = _T_6570[3]; // @[OneHot.scala 66:30:@3586.4]
  assign _T_6575 = _T_6570[4]; // @[OneHot.scala 66:30:@3587.4]
  assign _T_6576 = _T_6570[5]; // @[OneHot.scala 66:30:@3588.4]
  assign _T_6577 = _T_6570[6]; // @[OneHot.scala 66:30:@3589.4]
  assign _T_6578 = _T_6570[7]; // @[OneHot.scala 66:30:@3590.4]
  assign _T_6579 = _T_6570[8]; // @[OneHot.scala 66:30:@3591.4]
  assign _T_6580 = _T_6570[9]; // @[OneHot.scala 66:30:@3592.4]
  assign _T_6581 = _T_6570[10]; // @[OneHot.scala 66:30:@3593.4]
  assign _T_6582 = _T_6570[11]; // @[OneHot.scala 66:30:@3594.4]
  assign _T_6583 = _T_6570[12]; // @[OneHot.scala 66:30:@3595.4]
  assign _T_6584 = _T_6570[13]; // @[OneHot.scala 66:30:@3596.4]
  assign _T_6585 = _T_6570[14]; // @[OneHot.scala 66:30:@3597.4]
  assign _T_6586 = _T_6570[15]; // @[OneHot.scala 66:30:@3598.4]
  assign _T_6627 = _T_4217 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3616.4]
  assign _T_6628 = _T_4214 ? 16'h4000 : _T_6627; // @[Mux.scala 31:69:@3617.4]
  assign _T_6629 = _T_4211 ? 16'h2000 : _T_6628; // @[Mux.scala 31:69:@3618.4]
  assign _T_6630 = _T_4208 ? 16'h1000 : _T_6629; // @[Mux.scala 31:69:@3619.4]
  assign _T_6631 = _T_4205 ? 16'h800 : _T_6630; // @[Mux.scala 31:69:@3620.4]
  assign _T_6632 = _T_4202 ? 16'h400 : _T_6631; // @[Mux.scala 31:69:@3621.4]
  assign _T_6633 = _T_4199 ? 16'h200 : _T_6632; // @[Mux.scala 31:69:@3622.4]
  assign _T_6634 = _T_4196 ? 16'h100 : _T_6633; // @[Mux.scala 31:69:@3623.4]
  assign _T_6635 = _T_4193 ? 16'h80 : _T_6634; // @[Mux.scala 31:69:@3624.4]
  assign _T_6636 = _T_4238 ? 16'h40 : _T_6635; // @[Mux.scala 31:69:@3625.4]
  assign _T_6637 = _T_4235 ? 16'h20 : _T_6636; // @[Mux.scala 31:69:@3626.4]
  assign _T_6638 = _T_4232 ? 16'h10 : _T_6637; // @[Mux.scala 31:69:@3627.4]
  assign _T_6639 = _T_4229 ? 16'h8 : _T_6638; // @[Mux.scala 31:69:@3628.4]
  assign _T_6640 = _T_4226 ? 16'h4 : _T_6639; // @[Mux.scala 31:69:@3629.4]
  assign _T_6641 = _T_4223 ? 16'h2 : _T_6640; // @[Mux.scala 31:69:@3630.4]
  assign _T_6642 = _T_4220 ? 16'h1 : _T_6641; // @[Mux.scala 31:69:@3631.4]
  assign _T_6643 = _T_6642[0]; // @[OneHot.scala 66:30:@3632.4]
  assign _T_6644 = _T_6642[1]; // @[OneHot.scala 66:30:@3633.4]
  assign _T_6645 = _T_6642[2]; // @[OneHot.scala 66:30:@3634.4]
  assign _T_6646 = _T_6642[3]; // @[OneHot.scala 66:30:@3635.4]
  assign _T_6647 = _T_6642[4]; // @[OneHot.scala 66:30:@3636.4]
  assign _T_6648 = _T_6642[5]; // @[OneHot.scala 66:30:@3637.4]
  assign _T_6649 = _T_6642[6]; // @[OneHot.scala 66:30:@3638.4]
  assign _T_6650 = _T_6642[7]; // @[OneHot.scala 66:30:@3639.4]
  assign _T_6651 = _T_6642[8]; // @[OneHot.scala 66:30:@3640.4]
  assign _T_6652 = _T_6642[9]; // @[OneHot.scala 66:30:@3641.4]
  assign _T_6653 = _T_6642[10]; // @[OneHot.scala 66:30:@3642.4]
  assign _T_6654 = _T_6642[11]; // @[OneHot.scala 66:30:@3643.4]
  assign _T_6655 = _T_6642[12]; // @[OneHot.scala 66:30:@3644.4]
  assign _T_6656 = _T_6642[13]; // @[OneHot.scala 66:30:@3645.4]
  assign _T_6657 = _T_6642[14]; // @[OneHot.scala 66:30:@3646.4]
  assign _T_6658 = _T_6642[15]; // @[OneHot.scala 66:30:@3647.4]
  assign _T_6699 = _T_4220 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3665.4]
  assign _T_6700 = _T_4217 ? 16'h4000 : _T_6699; // @[Mux.scala 31:69:@3666.4]
  assign _T_6701 = _T_4214 ? 16'h2000 : _T_6700; // @[Mux.scala 31:69:@3667.4]
  assign _T_6702 = _T_4211 ? 16'h1000 : _T_6701; // @[Mux.scala 31:69:@3668.4]
  assign _T_6703 = _T_4208 ? 16'h800 : _T_6702; // @[Mux.scala 31:69:@3669.4]
  assign _T_6704 = _T_4205 ? 16'h400 : _T_6703; // @[Mux.scala 31:69:@3670.4]
  assign _T_6705 = _T_4202 ? 16'h200 : _T_6704; // @[Mux.scala 31:69:@3671.4]
  assign _T_6706 = _T_4199 ? 16'h100 : _T_6705; // @[Mux.scala 31:69:@3672.4]
  assign _T_6707 = _T_4196 ? 16'h80 : _T_6706; // @[Mux.scala 31:69:@3673.4]
  assign _T_6708 = _T_4193 ? 16'h40 : _T_6707; // @[Mux.scala 31:69:@3674.4]
  assign _T_6709 = _T_4238 ? 16'h20 : _T_6708; // @[Mux.scala 31:69:@3675.4]
  assign _T_6710 = _T_4235 ? 16'h10 : _T_6709; // @[Mux.scala 31:69:@3676.4]
  assign _T_6711 = _T_4232 ? 16'h8 : _T_6710; // @[Mux.scala 31:69:@3677.4]
  assign _T_6712 = _T_4229 ? 16'h4 : _T_6711; // @[Mux.scala 31:69:@3678.4]
  assign _T_6713 = _T_4226 ? 16'h2 : _T_6712; // @[Mux.scala 31:69:@3679.4]
  assign _T_6714 = _T_4223 ? 16'h1 : _T_6713; // @[Mux.scala 31:69:@3680.4]
  assign _T_6715 = _T_6714[0]; // @[OneHot.scala 66:30:@3681.4]
  assign _T_6716 = _T_6714[1]; // @[OneHot.scala 66:30:@3682.4]
  assign _T_6717 = _T_6714[2]; // @[OneHot.scala 66:30:@3683.4]
  assign _T_6718 = _T_6714[3]; // @[OneHot.scala 66:30:@3684.4]
  assign _T_6719 = _T_6714[4]; // @[OneHot.scala 66:30:@3685.4]
  assign _T_6720 = _T_6714[5]; // @[OneHot.scala 66:30:@3686.4]
  assign _T_6721 = _T_6714[6]; // @[OneHot.scala 66:30:@3687.4]
  assign _T_6722 = _T_6714[7]; // @[OneHot.scala 66:30:@3688.4]
  assign _T_6723 = _T_6714[8]; // @[OneHot.scala 66:30:@3689.4]
  assign _T_6724 = _T_6714[9]; // @[OneHot.scala 66:30:@3690.4]
  assign _T_6725 = _T_6714[10]; // @[OneHot.scala 66:30:@3691.4]
  assign _T_6726 = _T_6714[11]; // @[OneHot.scala 66:30:@3692.4]
  assign _T_6727 = _T_6714[12]; // @[OneHot.scala 66:30:@3693.4]
  assign _T_6728 = _T_6714[13]; // @[OneHot.scala 66:30:@3694.4]
  assign _T_6729 = _T_6714[14]; // @[OneHot.scala 66:30:@3695.4]
  assign _T_6730 = _T_6714[15]; // @[OneHot.scala 66:30:@3696.4]
  assign _T_6771 = _T_4223 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3714.4]
  assign _T_6772 = _T_4220 ? 16'h4000 : _T_6771; // @[Mux.scala 31:69:@3715.4]
  assign _T_6773 = _T_4217 ? 16'h2000 : _T_6772; // @[Mux.scala 31:69:@3716.4]
  assign _T_6774 = _T_4214 ? 16'h1000 : _T_6773; // @[Mux.scala 31:69:@3717.4]
  assign _T_6775 = _T_4211 ? 16'h800 : _T_6774; // @[Mux.scala 31:69:@3718.4]
  assign _T_6776 = _T_4208 ? 16'h400 : _T_6775; // @[Mux.scala 31:69:@3719.4]
  assign _T_6777 = _T_4205 ? 16'h200 : _T_6776; // @[Mux.scala 31:69:@3720.4]
  assign _T_6778 = _T_4202 ? 16'h100 : _T_6777; // @[Mux.scala 31:69:@3721.4]
  assign _T_6779 = _T_4199 ? 16'h80 : _T_6778; // @[Mux.scala 31:69:@3722.4]
  assign _T_6780 = _T_4196 ? 16'h40 : _T_6779; // @[Mux.scala 31:69:@3723.4]
  assign _T_6781 = _T_4193 ? 16'h20 : _T_6780; // @[Mux.scala 31:69:@3724.4]
  assign _T_6782 = _T_4238 ? 16'h10 : _T_6781; // @[Mux.scala 31:69:@3725.4]
  assign _T_6783 = _T_4235 ? 16'h8 : _T_6782; // @[Mux.scala 31:69:@3726.4]
  assign _T_6784 = _T_4232 ? 16'h4 : _T_6783; // @[Mux.scala 31:69:@3727.4]
  assign _T_6785 = _T_4229 ? 16'h2 : _T_6784; // @[Mux.scala 31:69:@3728.4]
  assign _T_6786 = _T_4226 ? 16'h1 : _T_6785; // @[Mux.scala 31:69:@3729.4]
  assign _T_6787 = _T_6786[0]; // @[OneHot.scala 66:30:@3730.4]
  assign _T_6788 = _T_6786[1]; // @[OneHot.scala 66:30:@3731.4]
  assign _T_6789 = _T_6786[2]; // @[OneHot.scala 66:30:@3732.4]
  assign _T_6790 = _T_6786[3]; // @[OneHot.scala 66:30:@3733.4]
  assign _T_6791 = _T_6786[4]; // @[OneHot.scala 66:30:@3734.4]
  assign _T_6792 = _T_6786[5]; // @[OneHot.scala 66:30:@3735.4]
  assign _T_6793 = _T_6786[6]; // @[OneHot.scala 66:30:@3736.4]
  assign _T_6794 = _T_6786[7]; // @[OneHot.scala 66:30:@3737.4]
  assign _T_6795 = _T_6786[8]; // @[OneHot.scala 66:30:@3738.4]
  assign _T_6796 = _T_6786[9]; // @[OneHot.scala 66:30:@3739.4]
  assign _T_6797 = _T_6786[10]; // @[OneHot.scala 66:30:@3740.4]
  assign _T_6798 = _T_6786[11]; // @[OneHot.scala 66:30:@3741.4]
  assign _T_6799 = _T_6786[12]; // @[OneHot.scala 66:30:@3742.4]
  assign _T_6800 = _T_6786[13]; // @[OneHot.scala 66:30:@3743.4]
  assign _T_6801 = _T_6786[14]; // @[OneHot.scala 66:30:@3744.4]
  assign _T_6802 = _T_6786[15]; // @[OneHot.scala 66:30:@3745.4]
  assign _T_6843 = _T_4226 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3763.4]
  assign _T_6844 = _T_4223 ? 16'h4000 : _T_6843; // @[Mux.scala 31:69:@3764.4]
  assign _T_6845 = _T_4220 ? 16'h2000 : _T_6844; // @[Mux.scala 31:69:@3765.4]
  assign _T_6846 = _T_4217 ? 16'h1000 : _T_6845; // @[Mux.scala 31:69:@3766.4]
  assign _T_6847 = _T_4214 ? 16'h800 : _T_6846; // @[Mux.scala 31:69:@3767.4]
  assign _T_6848 = _T_4211 ? 16'h400 : _T_6847; // @[Mux.scala 31:69:@3768.4]
  assign _T_6849 = _T_4208 ? 16'h200 : _T_6848; // @[Mux.scala 31:69:@3769.4]
  assign _T_6850 = _T_4205 ? 16'h100 : _T_6849; // @[Mux.scala 31:69:@3770.4]
  assign _T_6851 = _T_4202 ? 16'h80 : _T_6850; // @[Mux.scala 31:69:@3771.4]
  assign _T_6852 = _T_4199 ? 16'h40 : _T_6851; // @[Mux.scala 31:69:@3772.4]
  assign _T_6853 = _T_4196 ? 16'h20 : _T_6852; // @[Mux.scala 31:69:@3773.4]
  assign _T_6854 = _T_4193 ? 16'h10 : _T_6853; // @[Mux.scala 31:69:@3774.4]
  assign _T_6855 = _T_4238 ? 16'h8 : _T_6854; // @[Mux.scala 31:69:@3775.4]
  assign _T_6856 = _T_4235 ? 16'h4 : _T_6855; // @[Mux.scala 31:69:@3776.4]
  assign _T_6857 = _T_4232 ? 16'h2 : _T_6856; // @[Mux.scala 31:69:@3777.4]
  assign _T_6858 = _T_4229 ? 16'h1 : _T_6857; // @[Mux.scala 31:69:@3778.4]
  assign _T_6859 = _T_6858[0]; // @[OneHot.scala 66:30:@3779.4]
  assign _T_6860 = _T_6858[1]; // @[OneHot.scala 66:30:@3780.4]
  assign _T_6861 = _T_6858[2]; // @[OneHot.scala 66:30:@3781.4]
  assign _T_6862 = _T_6858[3]; // @[OneHot.scala 66:30:@3782.4]
  assign _T_6863 = _T_6858[4]; // @[OneHot.scala 66:30:@3783.4]
  assign _T_6864 = _T_6858[5]; // @[OneHot.scala 66:30:@3784.4]
  assign _T_6865 = _T_6858[6]; // @[OneHot.scala 66:30:@3785.4]
  assign _T_6866 = _T_6858[7]; // @[OneHot.scala 66:30:@3786.4]
  assign _T_6867 = _T_6858[8]; // @[OneHot.scala 66:30:@3787.4]
  assign _T_6868 = _T_6858[9]; // @[OneHot.scala 66:30:@3788.4]
  assign _T_6869 = _T_6858[10]; // @[OneHot.scala 66:30:@3789.4]
  assign _T_6870 = _T_6858[11]; // @[OneHot.scala 66:30:@3790.4]
  assign _T_6871 = _T_6858[12]; // @[OneHot.scala 66:30:@3791.4]
  assign _T_6872 = _T_6858[13]; // @[OneHot.scala 66:30:@3792.4]
  assign _T_6873 = _T_6858[14]; // @[OneHot.scala 66:30:@3793.4]
  assign _T_6874 = _T_6858[15]; // @[OneHot.scala 66:30:@3794.4]
  assign _T_6915 = _T_4229 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3812.4]
  assign _T_6916 = _T_4226 ? 16'h4000 : _T_6915; // @[Mux.scala 31:69:@3813.4]
  assign _T_6917 = _T_4223 ? 16'h2000 : _T_6916; // @[Mux.scala 31:69:@3814.4]
  assign _T_6918 = _T_4220 ? 16'h1000 : _T_6917; // @[Mux.scala 31:69:@3815.4]
  assign _T_6919 = _T_4217 ? 16'h800 : _T_6918; // @[Mux.scala 31:69:@3816.4]
  assign _T_6920 = _T_4214 ? 16'h400 : _T_6919; // @[Mux.scala 31:69:@3817.4]
  assign _T_6921 = _T_4211 ? 16'h200 : _T_6920; // @[Mux.scala 31:69:@3818.4]
  assign _T_6922 = _T_4208 ? 16'h100 : _T_6921; // @[Mux.scala 31:69:@3819.4]
  assign _T_6923 = _T_4205 ? 16'h80 : _T_6922; // @[Mux.scala 31:69:@3820.4]
  assign _T_6924 = _T_4202 ? 16'h40 : _T_6923; // @[Mux.scala 31:69:@3821.4]
  assign _T_6925 = _T_4199 ? 16'h20 : _T_6924; // @[Mux.scala 31:69:@3822.4]
  assign _T_6926 = _T_4196 ? 16'h10 : _T_6925; // @[Mux.scala 31:69:@3823.4]
  assign _T_6927 = _T_4193 ? 16'h8 : _T_6926; // @[Mux.scala 31:69:@3824.4]
  assign _T_6928 = _T_4238 ? 16'h4 : _T_6927; // @[Mux.scala 31:69:@3825.4]
  assign _T_6929 = _T_4235 ? 16'h2 : _T_6928; // @[Mux.scala 31:69:@3826.4]
  assign _T_6930 = _T_4232 ? 16'h1 : _T_6929; // @[Mux.scala 31:69:@3827.4]
  assign _T_6931 = _T_6930[0]; // @[OneHot.scala 66:30:@3828.4]
  assign _T_6932 = _T_6930[1]; // @[OneHot.scala 66:30:@3829.4]
  assign _T_6933 = _T_6930[2]; // @[OneHot.scala 66:30:@3830.4]
  assign _T_6934 = _T_6930[3]; // @[OneHot.scala 66:30:@3831.4]
  assign _T_6935 = _T_6930[4]; // @[OneHot.scala 66:30:@3832.4]
  assign _T_6936 = _T_6930[5]; // @[OneHot.scala 66:30:@3833.4]
  assign _T_6937 = _T_6930[6]; // @[OneHot.scala 66:30:@3834.4]
  assign _T_6938 = _T_6930[7]; // @[OneHot.scala 66:30:@3835.4]
  assign _T_6939 = _T_6930[8]; // @[OneHot.scala 66:30:@3836.4]
  assign _T_6940 = _T_6930[9]; // @[OneHot.scala 66:30:@3837.4]
  assign _T_6941 = _T_6930[10]; // @[OneHot.scala 66:30:@3838.4]
  assign _T_6942 = _T_6930[11]; // @[OneHot.scala 66:30:@3839.4]
  assign _T_6943 = _T_6930[12]; // @[OneHot.scala 66:30:@3840.4]
  assign _T_6944 = _T_6930[13]; // @[OneHot.scala 66:30:@3841.4]
  assign _T_6945 = _T_6930[14]; // @[OneHot.scala 66:30:@3842.4]
  assign _T_6946 = _T_6930[15]; // @[OneHot.scala 66:30:@3843.4]
  assign _T_6987 = _T_4232 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3861.4]
  assign _T_6988 = _T_4229 ? 16'h4000 : _T_6987; // @[Mux.scala 31:69:@3862.4]
  assign _T_6989 = _T_4226 ? 16'h2000 : _T_6988; // @[Mux.scala 31:69:@3863.4]
  assign _T_6990 = _T_4223 ? 16'h1000 : _T_6989; // @[Mux.scala 31:69:@3864.4]
  assign _T_6991 = _T_4220 ? 16'h800 : _T_6990; // @[Mux.scala 31:69:@3865.4]
  assign _T_6992 = _T_4217 ? 16'h400 : _T_6991; // @[Mux.scala 31:69:@3866.4]
  assign _T_6993 = _T_4214 ? 16'h200 : _T_6992; // @[Mux.scala 31:69:@3867.4]
  assign _T_6994 = _T_4211 ? 16'h100 : _T_6993; // @[Mux.scala 31:69:@3868.4]
  assign _T_6995 = _T_4208 ? 16'h80 : _T_6994; // @[Mux.scala 31:69:@3869.4]
  assign _T_6996 = _T_4205 ? 16'h40 : _T_6995; // @[Mux.scala 31:69:@3870.4]
  assign _T_6997 = _T_4202 ? 16'h20 : _T_6996; // @[Mux.scala 31:69:@3871.4]
  assign _T_6998 = _T_4199 ? 16'h10 : _T_6997; // @[Mux.scala 31:69:@3872.4]
  assign _T_6999 = _T_4196 ? 16'h8 : _T_6998; // @[Mux.scala 31:69:@3873.4]
  assign _T_7000 = _T_4193 ? 16'h4 : _T_6999; // @[Mux.scala 31:69:@3874.4]
  assign _T_7001 = _T_4238 ? 16'h2 : _T_7000; // @[Mux.scala 31:69:@3875.4]
  assign _T_7002 = _T_4235 ? 16'h1 : _T_7001; // @[Mux.scala 31:69:@3876.4]
  assign _T_7003 = _T_7002[0]; // @[OneHot.scala 66:30:@3877.4]
  assign _T_7004 = _T_7002[1]; // @[OneHot.scala 66:30:@3878.4]
  assign _T_7005 = _T_7002[2]; // @[OneHot.scala 66:30:@3879.4]
  assign _T_7006 = _T_7002[3]; // @[OneHot.scala 66:30:@3880.4]
  assign _T_7007 = _T_7002[4]; // @[OneHot.scala 66:30:@3881.4]
  assign _T_7008 = _T_7002[5]; // @[OneHot.scala 66:30:@3882.4]
  assign _T_7009 = _T_7002[6]; // @[OneHot.scala 66:30:@3883.4]
  assign _T_7010 = _T_7002[7]; // @[OneHot.scala 66:30:@3884.4]
  assign _T_7011 = _T_7002[8]; // @[OneHot.scala 66:30:@3885.4]
  assign _T_7012 = _T_7002[9]; // @[OneHot.scala 66:30:@3886.4]
  assign _T_7013 = _T_7002[10]; // @[OneHot.scala 66:30:@3887.4]
  assign _T_7014 = _T_7002[11]; // @[OneHot.scala 66:30:@3888.4]
  assign _T_7015 = _T_7002[12]; // @[OneHot.scala 66:30:@3889.4]
  assign _T_7016 = _T_7002[13]; // @[OneHot.scala 66:30:@3890.4]
  assign _T_7017 = _T_7002[14]; // @[OneHot.scala 66:30:@3891.4]
  assign _T_7018 = _T_7002[15]; // @[OneHot.scala 66:30:@3892.4]
  assign _T_7059 = _T_4235 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3910.4]
  assign _T_7060 = _T_4232 ? 16'h4000 : _T_7059; // @[Mux.scala 31:69:@3911.4]
  assign _T_7061 = _T_4229 ? 16'h2000 : _T_7060; // @[Mux.scala 31:69:@3912.4]
  assign _T_7062 = _T_4226 ? 16'h1000 : _T_7061; // @[Mux.scala 31:69:@3913.4]
  assign _T_7063 = _T_4223 ? 16'h800 : _T_7062; // @[Mux.scala 31:69:@3914.4]
  assign _T_7064 = _T_4220 ? 16'h400 : _T_7063; // @[Mux.scala 31:69:@3915.4]
  assign _T_7065 = _T_4217 ? 16'h200 : _T_7064; // @[Mux.scala 31:69:@3916.4]
  assign _T_7066 = _T_4214 ? 16'h100 : _T_7065; // @[Mux.scala 31:69:@3917.4]
  assign _T_7067 = _T_4211 ? 16'h80 : _T_7066; // @[Mux.scala 31:69:@3918.4]
  assign _T_7068 = _T_4208 ? 16'h40 : _T_7067; // @[Mux.scala 31:69:@3919.4]
  assign _T_7069 = _T_4205 ? 16'h20 : _T_7068; // @[Mux.scala 31:69:@3920.4]
  assign _T_7070 = _T_4202 ? 16'h10 : _T_7069; // @[Mux.scala 31:69:@3921.4]
  assign _T_7071 = _T_4199 ? 16'h8 : _T_7070; // @[Mux.scala 31:69:@3922.4]
  assign _T_7072 = _T_4196 ? 16'h4 : _T_7071; // @[Mux.scala 31:69:@3923.4]
  assign _T_7073 = _T_4193 ? 16'h2 : _T_7072; // @[Mux.scala 31:69:@3924.4]
  assign _T_7074 = _T_4238 ? 16'h1 : _T_7073; // @[Mux.scala 31:69:@3925.4]
  assign _T_7075 = _T_7074[0]; // @[OneHot.scala 66:30:@3926.4]
  assign _T_7076 = _T_7074[1]; // @[OneHot.scala 66:30:@3927.4]
  assign _T_7077 = _T_7074[2]; // @[OneHot.scala 66:30:@3928.4]
  assign _T_7078 = _T_7074[3]; // @[OneHot.scala 66:30:@3929.4]
  assign _T_7079 = _T_7074[4]; // @[OneHot.scala 66:30:@3930.4]
  assign _T_7080 = _T_7074[5]; // @[OneHot.scala 66:30:@3931.4]
  assign _T_7081 = _T_7074[6]; // @[OneHot.scala 66:30:@3932.4]
  assign _T_7082 = _T_7074[7]; // @[OneHot.scala 66:30:@3933.4]
  assign _T_7083 = _T_7074[8]; // @[OneHot.scala 66:30:@3934.4]
  assign _T_7084 = _T_7074[9]; // @[OneHot.scala 66:30:@3935.4]
  assign _T_7085 = _T_7074[10]; // @[OneHot.scala 66:30:@3936.4]
  assign _T_7086 = _T_7074[11]; // @[OneHot.scala 66:30:@3937.4]
  assign _T_7087 = _T_7074[12]; // @[OneHot.scala 66:30:@3938.4]
  assign _T_7088 = _T_7074[13]; // @[OneHot.scala 66:30:@3939.4]
  assign _T_7089 = _T_7074[14]; // @[OneHot.scala 66:30:@3940.4]
  assign _T_7090 = _T_7074[15]; // @[OneHot.scala 66:30:@3941.4]
  assign _T_7155 = {_T_6002,_T_6001,_T_6000,_T_5999,_T_5998,_T_5997,_T_5996,_T_5995}; // @[Mux.scala 19:72:@3965.4]
  assign _T_7163 = {_T_6010,_T_6009,_T_6008,_T_6007,_T_6006,_T_6005,_T_6004,_T_6003,_T_7155}; // @[Mux.scala 19:72:@3973.4]
  assign _T_7165 = _T_4265 ? _T_7163 : 16'h0; // @[Mux.scala 19:72:@3974.4]
  assign _T_7172 = {_T_6073,_T_6072,_T_6071,_T_6070,_T_6069,_T_6068,_T_6067,_T_6082}; // @[Mux.scala 19:72:@3981.4]
  assign _T_7180 = {_T_6081,_T_6080,_T_6079,_T_6078,_T_6077,_T_6076,_T_6075,_T_6074,_T_7172}; // @[Mux.scala 19:72:@3989.4]
  assign _T_7182 = _T_4266 ? _T_7180 : 16'h0; // @[Mux.scala 19:72:@3990.4]
  assign _T_7189 = {_T_6144,_T_6143,_T_6142,_T_6141,_T_6140,_T_6139,_T_6154,_T_6153}; // @[Mux.scala 19:72:@3997.4]
  assign _T_7197 = {_T_6152,_T_6151,_T_6150,_T_6149,_T_6148,_T_6147,_T_6146,_T_6145,_T_7189}; // @[Mux.scala 19:72:@4005.4]
  assign _T_7199 = _T_4267 ? _T_7197 : 16'h0; // @[Mux.scala 19:72:@4006.4]
  assign _T_7206 = {_T_6215,_T_6214,_T_6213,_T_6212,_T_6211,_T_6226,_T_6225,_T_6224}; // @[Mux.scala 19:72:@4013.4]
  assign _T_7214 = {_T_6223,_T_6222,_T_6221,_T_6220,_T_6219,_T_6218,_T_6217,_T_6216,_T_7206}; // @[Mux.scala 19:72:@4021.4]
  assign _T_7216 = _T_4268 ? _T_7214 : 16'h0; // @[Mux.scala 19:72:@4022.4]
  assign _T_7223 = {_T_6286,_T_6285,_T_6284,_T_6283,_T_6298,_T_6297,_T_6296,_T_6295}; // @[Mux.scala 19:72:@4029.4]
  assign _T_7231 = {_T_6294,_T_6293,_T_6292,_T_6291,_T_6290,_T_6289,_T_6288,_T_6287,_T_7223}; // @[Mux.scala 19:72:@4037.4]
  assign _T_7233 = _T_4269 ? _T_7231 : 16'h0; // @[Mux.scala 19:72:@4038.4]
  assign _T_7240 = {_T_6357,_T_6356,_T_6355,_T_6370,_T_6369,_T_6368,_T_6367,_T_6366}; // @[Mux.scala 19:72:@4045.4]
  assign _T_7248 = {_T_6365,_T_6364,_T_6363,_T_6362,_T_6361,_T_6360,_T_6359,_T_6358,_T_7240}; // @[Mux.scala 19:72:@4053.4]
  assign _T_7250 = _T_4270 ? _T_7248 : 16'h0; // @[Mux.scala 19:72:@4054.4]
  assign _T_7257 = {_T_6428,_T_6427,_T_6442,_T_6441,_T_6440,_T_6439,_T_6438,_T_6437}; // @[Mux.scala 19:72:@4061.4]
  assign _T_7265 = {_T_6436,_T_6435,_T_6434,_T_6433,_T_6432,_T_6431,_T_6430,_T_6429,_T_7257}; // @[Mux.scala 19:72:@4069.4]
  assign _T_7267 = _T_4271 ? _T_7265 : 16'h0; // @[Mux.scala 19:72:@4070.4]
  assign _T_7274 = {_T_6499,_T_6514,_T_6513,_T_6512,_T_6511,_T_6510,_T_6509,_T_6508}; // @[Mux.scala 19:72:@4077.4]
  assign _T_7282 = {_T_6507,_T_6506,_T_6505,_T_6504,_T_6503,_T_6502,_T_6501,_T_6500,_T_7274}; // @[Mux.scala 19:72:@4085.4]
  assign _T_7284 = _T_4272 ? _T_7282 : 16'h0; // @[Mux.scala 19:72:@4086.4]
  assign _T_7291 = {_T_6586,_T_6585,_T_6584,_T_6583,_T_6582,_T_6581,_T_6580,_T_6579}; // @[Mux.scala 19:72:@4093.4]
  assign _T_7299 = {_T_6578,_T_6577,_T_6576,_T_6575,_T_6574,_T_6573,_T_6572,_T_6571,_T_7291}; // @[Mux.scala 19:72:@4101.4]
  assign _T_7301 = _T_4273 ? _T_7299 : 16'h0; // @[Mux.scala 19:72:@4102.4]
  assign _T_7308 = {_T_6657,_T_6656,_T_6655,_T_6654,_T_6653,_T_6652,_T_6651,_T_6650}; // @[Mux.scala 19:72:@4109.4]
  assign _T_7316 = {_T_6649,_T_6648,_T_6647,_T_6646,_T_6645,_T_6644,_T_6643,_T_6658,_T_7308}; // @[Mux.scala 19:72:@4117.4]
  assign _T_7318 = _T_4274 ? _T_7316 : 16'h0; // @[Mux.scala 19:72:@4118.4]
  assign _T_7325 = {_T_6728,_T_6727,_T_6726,_T_6725,_T_6724,_T_6723,_T_6722,_T_6721}; // @[Mux.scala 19:72:@4125.4]
  assign _T_7333 = {_T_6720,_T_6719,_T_6718,_T_6717,_T_6716,_T_6715,_T_6730,_T_6729,_T_7325}; // @[Mux.scala 19:72:@4133.4]
  assign _T_7335 = _T_4275 ? _T_7333 : 16'h0; // @[Mux.scala 19:72:@4134.4]
  assign _T_7342 = {_T_6799,_T_6798,_T_6797,_T_6796,_T_6795,_T_6794,_T_6793,_T_6792}; // @[Mux.scala 19:72:@4141.4]
  assign _T_7350 = {_T_6791,_T_6790,_T_6789,_T_6788,_T_6787,_T_6802,_T_6801,_T_6800,_T_7342}; // @[Mux.scala 19:72:@4149.4]
  assign _T_7352 = _T_4276 ? _T_7350 : 16'h0; // @[Mux.scala 19:72:@4150.4]
  assign _T_7359 = {_T_6870,_T_6869,_T_6868,_T_6867,_T_6866,_T_6865,_T_6864,_T_6863}; // @[Mux.scala 19:72:@4157.4]
  assign _T_7367 = {_T_6862,_T_6861,_T_6860,_T_6859,_T_6874,_T_6873,_T_6872,_T_6871,_T_7359}; // @[Mux.scala 19:72:@4165.4]
  assign _T_7369 = _T_4277 ? _T_7367 : 16'h0; // @[Mux.scala 19:72:@4166.4]
  assign _T_7376 = {_T_6941,_T_6940,_T_6939,_T_6938,_T_6937,_T_6936,_T_6935,_T_6934}; // @[Mux.scala 19:72:@4173.4]
  assign _T_7384 = {_T_6933,_T_6932,_T_6931,_T_6946,_T_6945,_T_6944,_T_6943,_T_6942,_T_7376}; // @[Mux.scala 19:72:@4181.4]
  assign _T_7386 = _T_4278 ? _T_7384 : 16'h0; // @[Mux.scala 19:72:@4182.4]
  assign _T_7393 = {_T_7012,_T_7011,_T_7010,_T_7009,_T_7008,_T_7007,_T_7006,_T_7005}; // @[Mux.scala 19:72:@4189.4]
  assign _T_7401 = {_T_7004,_T_7003,_T_7018,_T_7017,_T_7016,_T_7015,_T_7014,_T_7013,_T_7393}; // @[Mux.scala 19:72:@4197.4]
  assign _T_7403 = _T_4279 ? _T_7401 : 16'h0; // @[Mux.scala 19:72:@4198.4]
  assign _T_7410 = {_T_7083,_T_7082,_T_7081,_T_7080,_T_7079,_T_7078,_T_7077,_T_7076}; // @[Mux.scala 19:72:@4205.4]
  assign _T_7418 = {_T_7075,_T_7090,_T_7089,_T_7088,_T_7087,_T_7086,_T_7085,_T_7084,_T_7410}; // @[Mux.scala 19:72:@4213.4]
  assign _T_7420 = _T_4280 ? _T_7418 : 16'h0; // @[Mux.scala 19:72:@4214.4]
  assign _T_7421 = _T_7165 | _T_7182; // @[Mux.scala 19:72:@4215.4]
  assign _T_7422 = _T_7421 | _T_7199; // @[Mux.scala 19:72:@4216.4]
  assign _T_7423 = _T_7422 | _T_7216; // @[Mux.scala 19:72:@4217.4]
  assign _T_7424 = _T_7423 | _T_7233; // @[Mux.scala 19:72:@4218.4]
  assign _T_7425 = _T_7424 | _T_7250; // @[Mux.scala 19:72:@4219.4]
  assign _T_7426 = _T_7425 | _T_7267; // @[Mux.scala 19:72:@4220.4]
  assign _T_7427 = _T_7426 | _T_7284; // @[Mux.scala 19:72:@4221.4]
  assign _T_7428 = _T_7427 | _T_7301; // @[Mux.scala 19:72:@4222.4]
  assign _T_7429 = _T_7428 | _T_7318; // @[Mux.scala 19:72:@4223.4]
  assign _T_7430 = _T_7429 | _T_7335; // @[Mux.scala 19:72:@4224.4]
  assign _T_7431 = _T_7430 | _T_7352; // @[Mux.scala 19:72:@4225.4]
  assign _T_7432 = _T_7431 | _T_7369; // @[Mux.scala 19:72:@4226.4]
  assign _T_7433 = _T_7432 | _T_7386; // @[Mux.scala 19:72:@4227.4]
  assign _T_7434 = _T_7433 | _T_7403; // @[Mux.scala 19:72:@4228.4]
  assign _T_7435 = _T_7434 | _T_7420; // @[Mux.scala 19:72:@4229.4]
  assign inputDataPriorityPorts_0_0 = _T_7435[0]; // @[Mux.scala 19:72:@4233.4]
  assign inputDataPriorityPorts_0_1 = _T_7435[1]; // @[Mux.scala 19:72:@4235.4]
  assign inputDataPriorityPorts_0_2 = _T_7435[2]; // @[Mux.scala 19:72:@4237.4]
  assign inputDataPriorityPorts_0_3 = _T_7435[3]; // @[Mux.scala 19:72:@4239.4]
  assign inputDataPriorityPorts_0_4 = _T_7435[4]; // @[Mux.scala 19:72:@4241.4]
  assign inputDataPriorityPorts_0_5 = _T_7435[5]; // @[Mux.scala 19:72:@4243.4]
  assign inputDataPriorityPorts_0_6 = _T_7435[6]; // @[Mux.scala 19:72:@4245.4]
  assign inputDataPriorityPorts_0_7 = _T_7435[7]; // @[Mux.scala 19:72:@4247.4]
  assign inputDataPriorityPorts_0_8 = _T_7435[8]; // @[Mux.scala 19:72:@4249.4]
  assign inputDataPriorityPorts_0_9 = _T_7435[9]; // @[Mux.scala 19:72:@4251.4]
  assign inputDataPriorityPorts_0_10 = _T_7435[10]; // @[Mux.scala 19:72:@4253.4]
  assign inputDataPriorityPorts_0_11 = _T_7435[11]; // @[Mux.scala 19:72:@4255.4]
  assign inputDataPriorityPorts_0_12 = _T_7435[12]; // @[Mux.scala 19:72:@4257.4]
  assign inputDataPriorityPorts_0_13 = _T_7435[13]; // @[Mux.scala 19:72:@4259.4]
  assign inputDataPriorityPorts_0_14 = _T_7435[14]; // @[Mux.scala 19:72:@4261.4]
  assign inputDataPriorityPorts_0_15 = _T_7435[15]; // @[Mux.scala 19:72:@4263.4]
  assign _T_7581 = inputAddrPriorityPorts_0_0 & _T_4122; // @[StoreQueue.scala 209:52:@4287.6]
  assign _T_7582 = _T_7581 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4288.6]
  assign _GEN_992 = _T_7582 ? io_addressFromStorePorts_0 : addrQ_0; // @[StoreQueue.scala 210:40:@4292.6]
  assign _GEN_993 = _T_7582 ? 1'h1 : addrKnown_0; // @[StoreQueue.scala 210:40:@4292.6]
  assign _T_7598 = inputDataPriorityPorts_0_0 & _T_4192; // @[StoreQueue.scala 215:52:@4297.6]
  assign _T_7599 = _T_7598 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4298.6]
  assign _GEN_994 = _T_7599 ? io_dataFromStorePorts_0 : dataQ_0; // @[StoreQueue.scala 216:40:@4302.6]
  assign _GEN_995 = _T_7599 ? 1'h1 : dataKnown_0; // @[StoreQueue.scala 216:40:@4302.6]
  assign _GEN_996 = initBits_0 ? 1'h0 : _GEN_993; // @[StoreQueue.scala 204:35:@4281.4]
  assign _GEN_997 = initBits_0 ? 1'h0 : _GEN_995; // @[StoreQueue.scala 204:35:@4281.4]
  assign _GEN_998 = initBits_0 ? addrQ_0 : _GEN_992; // @[StoreQueue.scala 204:35:@4281.4]
  assign _GEN_999 = initBits_0 ? dataQ_0 : _GEN_994; // @[StoreQueue.scala 204:35:@4281.4]
  assign _T_7617 = inputAddrPriorityPorts_0_1 & _T_4125; // @[StoreQueue.scala 209:52:@4313.6]
  assign _T_7618 = _T_7617 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4314.6]
  assign _GEN_1000 = _T_7618 ? io_addressFromStorePorts_0 : addrQ_1; // @[StoreQueue.scala 210:40:@4318.6]
  assign _GEN_1001 = _T_7618 ? 1'h1 : addrKnown_1; // @[StoreQueue.scala 210:40:@4318.6]
  assign _T_7634 = inputDataPriorityPorts_0_1 & _T_4195; // @[StoreQueue.scala 215:52:@4323.6]
  assign _T_7635 = _T_7634 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4324.6]
  assign _GEN_1002 = _T_7635 ? io_dataFromStorePorts_0 : dataQ_1; // @[StoreQueue.scala 216:40:@4328.6]
  assign _GEN_1003 = _T_7635 ? 1'h1 : dataKnown_1; // @[StoreQueue.scala 216:40:@4328.6]
  assign _GEN_1004 = initBits_1 ? 1'h0 : _GEN_1001; // @[StoreQueue.scala 204:35:@4307.4]
  assign _GEN_1005 = initBits_1 ? 1'h0 : _GEN_1003; // @[StoreQueue.scala 204:35:@4307.4]
  assign _GEN_1006 = initBits_1 ? addrQ_1 : _GEN_1000; // @[StoreQueue.scala 204:35:@4307.4]
  assign _GEN_1007 = initBits_1 ? dataQ_1 : _GEN_1002; // @[StoreQueue.scala 204:35:@4307.4]
  assign _T_7653 = inputAddrPriorityPorts_0_2 & _T_4128; // @[StoreQueue.scala 209:52:@4339.6]
  assign _T_7654 = _T_7653 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4340.6]
  assign _GEN_1008 = _T_7654 ? io_addressFromStorePorts_0 : addrQ_2; // @[StoreQueue.scala 210:40:@4344.6]
  assign _GEN_1009 = _T_7654 ? 1'h1 : addrKnown_2; // @[StoreQueue.scala 210:40:@4344.6]
  assign _T_7670 = inputDataPriorityPorts_0_2 & _T_4198; // @[StoreQueue.scala 215:52:@4349.6]
  assign _T_7671 = _T_7670 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4350.6]
  assign _GEN_1010 = _T_7671 ? io_dataFromStorePorts_0 : dataQ_2; // @[StoreQueue.scala 216:40:@4354.6]
  assign _GEN_1011 = _T_7671 ? 1'h1 : dataKnown_2; // @[StoreQueue.scala 216:40:@4354.6]
  assign _GEN_1012 = initBits_2 ? 1'h0 : _GEN_1009; // @[StoreQueue.scala 204:35:@4333.4]
  assign _GEN_1013 = initBits_2 ? 1'h0 : _GEN_1011; // @[StoreQueue.scala 204:35:@4333.4]
  assign _GEN_1014 = initBits_2 ? addrQ_2 : _GEN_1008; // @[StoreQueue.scala 204:35:@4333.4]
  assign _GEN_1015 = initBits_2 ? dataQ_2 : _GEN_1010; // @[StoreQueue.scala 204:35:@4333.4]
  assign _T_7689 = inputAddrPriorityPorts_0_3 & _T_4131; // @[StoreQueue.scala 209:52:@4365.6]
  assign _T_7690 = _T_7689 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4366.6]
  assign _GEN_1016 = _T_7690 ? io_addressFromStorePorts_0 : addrQ_3; // @[StoreQueue.scala 210:40:@4370.6]
  assign _GEN_1017 = _T_7690 ? 1'h1 : addrKnown_3; // @[StoreQueue.scala 210:40:@4370.6]
  assign _T_7706 = inputDataPriorityPorts_0_3 & _T_4201; // @[StoreQueue.scala 215:52:@4375.6]
  assign _T_7707 = _T_7706 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4376.6]
  assign _GEN_1018 = _T_7707 ? io_dataFromStorePorts_0 : dataQ_3; // @[StoreQueue.scala 216:40:@4380.6]
  assign _GEN_1019 = _T_7707 ? 1'h1 : dataKnown_3; // @[StoreQueue.scala 216:40:@4380.6]
  assign _GEN_1020 = initBits_3 ? 1'h0 : _GEN_1017; // @[StoreQueue.scala 204:35:@4359.4]
  assign _GEN_1021 = initBits_3 ? 1'h0 : _GEN_1019; // @[StoreQueue.scala 204:35:@4359.4]
  assign _GEN_1022 = initBits_3 ? addrQ_3 : _GEN_1016; // @[StoreQueue.scala 204:35:@4359.4]
  assign _GEN_1023 = initBits_3 ? dataQ_3 : _GEN_1018; // @[StoreQueue.scala 204:35:@4359.4]
  assign _T_7725 = inputAddrPriorityPorts_0_4 & _T_4134; // @[StoreQueue.scala 209:52:@4391.6]
  assign _T_7726 = _T_7725 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4392.6]
  assign _GEN_1024 = _T_7726 ? io_addressFromStorePorts_0 : addrQ_4; // @[StoreQueue.scala 210:40:@4396.6]
  assign _GEN_1025 = _T_7726 ? 1'h1 : addrKnown_4; // @[StoreQueue.scala 210:40:@4396.6]
  assign _T_7742 = inputDataPriorityPorts_0_4 & _T_4204; // @[StoreQueue.scala 215:52:@4401.6]
  assign _T_7743 = _T_7742 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4402.6]
  assign _GEN_1026 = _T_7743 ? io_dataFromStorePorts_0 : dataQ_4; // @[StoreQueue.scala 216:40:@4406.6]
  assign _GEN_1027 = _T_7743 ? 1'h1 : dataKnown_4; // @[StoreQueue.scala 216:40:@4406.6]
  assign _GEN_1028 = initBits_4 ? 1'h0 : _GEN_1025; // @[StoreQueue.scala 204:35:@4385.4]
  assign _GEN_1029 = initBits_4 ? 1'h0 : _GEN_1027; // @[StoreQueue.scala 204:35:@4385.4]
  assign _GEN_1030 = initBits_4 ? addrQ_4 : _GEN_1024; // @[StoreQueue.scala 204:35:@4385.4]
  assign _GEN_1031 = initBits_4 ? dataQ_4 : _GEN_1026; // @[StoreQueue.scala 204:35:@4385.4]
  assign _T_7761 = inputAddrPriorityPorts_0_5 & _T_4137; // @[StoreQueue.scala 209:52:@4417.6]
  assign _T_7762 = _T_7761 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4418.6]
  assign _GEN_1032 = _T_7762 ? io_addressFromStorePorts_0 : addrQ_5; // @[StoreQueue.scala 210:40:@4422.6]
  assign _GEN_1033 = _T_7762 ? 1'h1 : addrKnown_5; // @[StoreQueue.scala 210:40:@4422.6]
  assign _T_7778 = inputDataPriorityPorts_0_5 & _T_4207; // @[StoreQueue.scala 215:52:@4427.6]
  assign _T_7779 = _T_7778 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4428.6]
  assign _GEN_1034 = _T_7779 ? io_dataFromStorePorts_0 : dataQ_5; // @[StoreQueue.scala 216:40:@4432.6]
  assign _GEN_1035 = _T_7779 ? 1'h1 : dataKnown_5; // @[StoreQueue.scala 216:40:@4432.6]
  assign _GEN_1036 = initBits_5 ? 1'h0 : _GEN_1033; // @[StoreQueue.scala 204:35:@4411.4]
  assign _GEN_1037 = initBits_5 ? 1'h0 : _GEN_1035; // @[StoreQueue.scala 204:35:@4411.4]
  assign _GEN_1038 = initBits_5 ? addrQ_5 : _GEN_1032; // @[StoreQueue.scala 204:35:@4411.4]
  assign _GEN_1039 = initBits_5 ? dataQ_5 : _GEN_1034; // @[StoreQueue.scala 204:35:@4411.4]
  assign _T_7797 = inputAddrPriorityPorts_0_6 & _T_4140; // @[StoreQueue.scala 209:52:@4443.6]
  assign _T_7798 = _T_7797 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4444.6]
  assign _GEN_1040 = _T_7798 ? io_addressFromStorePorts_0 : addrQ_6; // @[StoreQueue.scala 210:40:@4448.6]
  assign _GEN_1041 = _T_7798 ? 1'h1 : addrKnown_6; // @[StoreQueue.scala 210:40:@4448.6]
  assign _T_7814 = inputDataPriorityPorts_0_6 & _T_4210; // @[StoreQueue.scala 215:52:@4453.6]
  assign _T_7815 = _T_7814 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4454.6]
  assign _GEN_1042 = _T_7815 ? io_dataFromStorePorts_0 : dataQ_6; // @[StoreQueue.scala 216:40:@4458.6]
  assign _GEN_1043 = _T_7815 ? 1'h1 : dataKnown_6; // @[StoreQueue.scala 216:40:@4458.6]
  assign _GEN_1044 = initBits_6 ? 1'h0 : _GEN_1041; // @[StoreQueue.scala 204:35:@4437.4]
  assign _GEN_1045 = initBits_6 ? 1'h0 : _GEN_1043; // @[StoreQueue.scala 204:35:@4437.4]
  assign _GEN_1046 = initBits_6 ? addrQ_6 : _GEN_1040; // @[StoreQueue.scala 204:35:@4437.4]
  assign _GEN_1047 = initBits_6 ? dataQ_6 : _GEN_1042; // @[StoreQueue.scala 204:35:@4437.4]
  assign _T_7833 = inputAddrPriorityPorts_0_7 & _T_4143; // @[StoreQueue.scala 209:52:@4469.6]
  assign _T_7834 = _T_7833 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4470.6]
  assign _GEN_1048 = _T_7834 ? io_addressFromStorePorts_0 : addrQ_7; // @[StoreQueue.scala 210:40:@4474.6]
  assign _GEN_1049 = _T_7834 ? 1'h1 : addrKnown_7; // @[StoreQueue.scala 210:40:@4474.6]
  assign _T_7850 = inputDataPriorityPorts_0_7 & _T_4213; // @[StoreQueue.scala 215:52:@4479.6]
  assign _T_7851 = _T_7850 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4480.6]
  assign _GEN_1050 = _T_7851 ? io_dataFromStorePorts_0 : dataQ_7; // @[StoreQueue.scala 216:40:@4484.6]
  assign _GEN_1051 = _T_7851 ? 1'h1 : dataKnown_7; // @[StoreQueue.scala 216:40:@4484.6]
  assign _GEN_1052 = initBits_7 ? 1'h0 : _GEN_1049; // @[StoreQueue.scala 204:35:@4463.4]
  assign _GEN_1053 = initBits_7 ? 1'h0 : _GEN_1051; // @[StoreQueue.scala 204:35:@4463.4]
  assign _GEN_1054 = initBits_7 ? addrQ_7 : _GEN_1048; // @[StoreQueue.scala 204:35:@4463.4]
  assign _GEN_1055 = initBits_7 ? dataQ_7 : _GEN_1050; // @[StoreQueue.scala 204:35:@4463.4]
  assign _T_7869 = inputAddrPriorityPorts_0_8 & _T_4146; // @[StoreQueue.scala 209:52:@4495.6]
  assign _T_7870 = _T_7869 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4496.6]
  assign _GEN_1056 = _T_7870 ? io_addressFromStorePorts_0 : addrQ_8; // @[StoreQueue.scala 210:40:@4500.6]
  assign _GEN_1057 = _T_7870 ? 1'h1 : addrKnown_8; // @[StoreQueue.scala 210:40:@4500.6]
  assign _T_7886 = inputDataPriorityPorts_0_8 & _T_4216; // @[StoreQueue.scala 215:52:@4505.6]
  assign _T_7887 = _T_7886 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4506.6]
  assign _GEN_1058 = _T_7887 ? io_dataFromStorePorts_0 : dataQ_8; // @[StoreQueue.scala 216:40:@4510.6]
  assign _GEN_1059 = _T_7887 ? 1'h1 : dataKnown_8; // @[StoreQueue.scala 216:40:@4510.6]
  assign _GEN_1060 = initBits_8 ? 1'h0 : _GEN_1057; // @[StoreQueue.scala 204:35:@4489.4]
  assign _GEN_1061 = initBits_8 ? 1'h0 : _GEN_1059; // @[StoreQueue.scala 204:35:@4489.4]
  assign _GEN_1062 = initBits_8 ? addrQ_8 : _GEN_1056; // @[StoreQueue.scala 204:35:@4489.4]
  assign _GEN_1063 = initBits_8 ? dataQ_8 : _GEN_1058; // @[StoreQueue.scala 204:35:@4489.4]
  assign _T_7905 = inputAddrPriorityPorts_0_9 & _T_4149; // @[StoreQueue.scala 209:52:@4521.6]
  assign _T_7906 = _T_7905 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4522.6]
  assign _GEN_1064 = _T_7906 ? io_addressFromStorePorts_0 : addrQ_9; // @[StoreQueue.scala 210:40:@4526.6]
  assign _GEN_1065 = _T_7906 ? 1'h1 : addrKnown_9; // @[StoreQueue.scala 210:40:@4526.6]
  assign _T_7922 = inputDataPriorityPorts_0_9 & _T_4219; // @[StoreQueue.scala 215:52:@4531.6]
  assign _T_7923 = _T_7922 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4532.6]
  assign _GEN_1066 = _T_7923 ? io_dataFromStorePorts_0 : dataQ_9; // @[StoreQueue.scala 216:40:@4536.6]
  assign _GEN_1067 = _T_7923 ? 1'h1 : dataKnown_9; // @[StoreQueue.scala 216:40:@4536.6]
  assign _GEN_1068 = initBits_9 ? 1'h0 : _GEN_1065; // @[StoreQueue.scala 204:35:@4515.4]
  assign _GEN_1069 = initBits_9 ? 1'h0 : _GEN_1067; // @[StoreQueue.scala 204:35:@4515.4]
  assign _GEN_1070 = initBits_9 ? addrQ_9 : _GEN_1064; // @[StoreQueue.scala 204:35:@4515.4]
  assign _GEN_1071 = initBits_9 ? dataQ_9 : _GEN_1066; // @[StoreQueue.scala 204:35:@4515.4]
  assign _T_7941 = inputAddrPriorityPorts_0_10 & _T_4152; // @[StoreQueue.scala 209:52:@4547.6]
  assign _T_7942 = _T_7941 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4548.6]
  assign _GEN_1072 = _T_7942 ? io_addressFromStorePorts_0 : addrQ_10; // @[StoreQueue.scala 210:40:@4552.6]
  assign _GEN_1073 = _T_7942 ? 1'h1 : addrKnown_10; // @[StoreQueue.scala 210:40:@4552.6]
  assign _T_7958 = inputDataPriorityPorts_0_10 & _T_4222; // @[StoreQueue.scala 215:52:@4557.6]
  assign _T_7959 = _T_7958 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4558.6]
  assign _GEN_1074 = _T_7959 ? io_dataFromStorePorts_0 : dataQ_10; // @[StoreQueue.scala 216:40:@4562.6]
  assign _GEN_1075 = _T_7959 ? 1'h1 : dataKnown_10; // @[StoreQueue.scala 216:40:@4562.6]
  assign _GEN_1076 = initBits_10 ? 1'h0 : _GEN_1073; // @[StoreQueue.scala 204:35:@4541.4]
  assign _GEN_1077 = initBits_10 ? 1'h0 : _GEN_1075; // @[StoreQueue.scala 204:35:@4541.4]
  assign _GEN_1078 = initBits_10 ? addrQ_10 : _GEN_1072; // @[StoreQueue.scala 204:35:@4541.4]
  assign _GEN_1079 = initBits_10 ? dataQ_10 : _GEN_1074; // @[StoreQueue.scala 204:35:@4541.4]
  assign _T_7977 = inputAddrPriorityPorts_0_11 & _T_4155; // @[StoreQueue.scala 209:52:@4573.6]
  assign _T_7978 = _T_7977 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4574.6]
  assign _GEN_1080 = _T_7978 ? io_addressFromStorePorts_0 : addrQ_11; // @[StoreQueue.scala 210:40:@4578.6]
  assign _GEN_1081 = _T_7978 ? 1'h1 : addrKnown_11; // @[StoreQueue.scala 210:40:@4578.6]
  assign _T_7994 = inputDataPriorityPorts_0_11 & _T_4225; // @[StoreQueue.scala 215:52:@4583.6]
  assign _T_7995 = _T_7994 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4584.6]
  assign _GEN_1082 = _T_7995 ? io_dataFromStorePorts_0 : dataQ_11; // @[StoreQueue.scala 216:40:@4588.6]
  assign _GEN_1083 = _T_7995 ? 1'h1 : dataKnown_11; // @[StoreQueue.scala 216:40:@4588.6]
  assign _GEN_1084 = initBits_11 ? 1'h0 : _GEN_1081; // @[StoreQueue.scala 204:35:@4567.4]
  assign _GEN_1085 = initBits_11 ? 1'h0 : _GEN_1083; // @[StoreQueue.scala 204:35:@4567.4]
  assign _GEN_1086 = initBits_11 ? addrQ_11 : _GEN_1080; // @[StoreQueue.scala 204:35:@4567.4]
  assign _GEN_1087 = initBits_11 ? dataQ_11 : _GEN_1082; // @[StoreQueue.scala 204:35:@4567.4]
  assign _T_8013 = inputAddrPriorityPorts_0_12 & _T_4158; // @[StoreQueue.scala 209:52:@4599.6]
  assign _T_8014 = _T_8013 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4600.6]
  assign _GEN_1088 = _T_8014 ? io_addressFromStorePorts_0 : addrQ_12; // @[StoreQueue.scala 210:40:@4604.6]
  assign _GEN_1089 = _T_8014 ? 1'h1 : addrKnown_12; // @[StoreQueue.scala 210:40:@4604.6]
  assign _T_8030 = inputDataPriorityPorts_0_12 & _T_4228; // @[StoreQueue.scala 215:52:@4609.6]
  assign _T_8031 = _T_8030 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4610.6]
  assign _GEN_1090 = _T_8031 ? io_dataFromStorePorts_0 : dataQ_12; // @[StoreQueue.scala 216:40:@4614.6]
  assign _GEN_1091 = _T_8031 ? 1'h1 : dataKnown_12; // @[StoreQueue.scala 216:40:@4614.6]
  assign _GEN_1092 = initBits_12 ? 1'h0 : _GEN_1089; // @[StoreQueue.scala 204:35:@4593.4]
  assign _GEN_1093 = initBits_12 ? 1'h0 : _GEN_1091; // @[StoreQueue.scala 204:35:@4593.4]
  assign _GEN_1094 = initBits_12 ? addrQ_12 : _GEN_1088; // @[StoreQueue.scala 204:35:@4593.4]
  assign _GEN_1095 = initBits_12 ? dataQ_12 : _GEN_1090; // @[StoreQueue.scala 204:35:@4593.4]
  assign _T_8049 = inputAddrPriorityPorts_0_13 & _T_4161; // @[StoreQueue.scala 209:52:@4625.6]
  assign _T_8050 = _T_8049 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4626.6]
  assign _GEN_1096 = _T_8050 ? io_addressFromStorePorts_0 : addrQ_13; // @[StoreQueue.scala 210:40:@4630.6]
  assign _GEN_1097 = _T_8050 ? 1'h1 : addrKnown_13; // @[StoreQueue.scala 210:40:@4630.6]
  assign _T_8066 = inputDataPriorityPorts_0_13 & _T_4231; // @[StoreQueue.scala 215:52:@4635.6]
  assign _T_8067 = _T_8066 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4636.6]
  assign _GEN_1098 = _T_8067 ? io_dataFromStorePorts_0 : dataQ_13; // @[StoreQueue.scala 216:40:@4640.6]
  assign _GEN_1099 = _T_8067 ? 1'h1 : dataKnown_13; // @[StoreQueue.scala 216:40:@4640.6]
  assign _GEN_1100 = initBits_13 ? 1'h0 : _GEN_1097; // @[StoreQueue.scala 204:35:@4619.4]
  assign _GEN_1101 = initBits_13 ? 1'h0 : _GEN_1099; // @[StoreQueue.scala 204:35:@4619.4]
  assign _GEN_1102 = initBits_13 ? addrQ_13 : _GEN_1096; // @[StoreQueue.scala 204:35:@4619.4]
  assign _GEN_1103 = initBits_13 ? dataQ_13 : _GEN_1098; // @[StoreQueue.scala 204:35:@4619.4]
  assign _T_8085 = inputAddrPriorityPorts_0_14 & _T_4164; // @[StoreQueue.scala 209:52:@4651.6]
  assign _T_8086 = _T_8085 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4652.6]
  assign _GEN_1104 = _T_8086 ? io_addressFromStorePorts_0 : addrQ_14; // @[StoreQueue.scala 210:40:@4656.6]
  assign _GEN_1105 = _T_8086 ? 1'h1 : addrKnown_14; // @[StoreQueue.scala 210:40:@4656.6]
  assign _T_8102 = inputDataPriorityPorts_0_14 & _T_4234; // @[StoreQueue.scala 215:52:@4661.6]
  assign _T_8103 = _T_8102 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4662.6]
  assign _GEN_1106 = _T_8103 ? io_dataFromStorePorts_0 : dataQ_14; // @[StoreQueue.scala 216:40:@4666.6]
  assign _GEN_1107 = _T_8103 ? 1'h1 : dataKnown_14; // @[StoreQueue.scala 216:40:@4666.6]
  assign _GEN_1108 = initBits_14 ? 1'h0 : _GEN_1105; // @[StoreQueue.scala 204:35:@4645.4]
  assign _GEN_1109 = initBits_14 ? 1'h0 : _GEN_1107; // @[StoreQueue.scala 204:35:@4645.4]
  assign _GEN_1110 = initBits_14 ? addrQ_14 : _GEN_1104; // @[StoreQueue.scala 204:35:@4645.4]
  assign _GEN_1111 = initBits_14 ? dataQ_14 : _GEN_1106; // @[StoreQueue.scala 204:35:@4645.4]
  assign _T_8121 = inputAddrPriorityPorts_0_15 & _T_4167; // @[StoreQueue.scala 209:52:@4677.6]
  assign _T_8122 = _T_8121 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4678.6]
  assign _GEN_1112 = _T_8122 ? io_addressFromStorePorts_0 : addrQ_15; // @[StoreQueue.scala 210:40:@4682.6]
  assign _GEN_1113 = _T_8122 ? 1'h1 : addrKnown_15; // @[StoreQueue.scala 210:40:@4682.6]
  assign _T_8138 = inputDataPriorityPorts_0_15 & _T_4237; // @[StoreQueue.scala 215:52:@4687.6]
  assign _T_8139 = _T_8138 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4688.6]
  assign _GEN_1114 = _T_8139 ? io_dataFromStorePorts_0 : dataQ_15; // @[StoreQueue.scala 216:40:@4692.6]
  assign _GEN_1115 = _T_8139 ? 1'h1 : dataKnown_15; // @[StoreQueue.scala 216:40:@4692.6]
  assign _GEN_1116 = initBits_15 ? 1'h0 : _GEN_1113; // @[StoreQueue.scala 204:35:@4671.4]
  assign _GEN_1117 = initBits_15 ? 1'h0 : _GEN_1115; // @[StoreQueue.scala 204:35:@4671.4]
  assign _GEN_1118 = initBits_15 ? addrQ_15 : _GEN_1112; // @[StoreQueue.scala 204:35:@4671.4]
  assign _GEN_1119 = initBits_15 ? dataQ_15 : _GEN_1114; // @[StoreQueue.scala 204:35:@4671.4]
  assign _T_8153 = storeRequest & io_memIsReadyForStores; // @[StoreQueue.scala 229:23:@4697.4]
  assign _T_8156 = head + 4'h1; // @[util.scala 10:8:@4699.6]
  assign _GEN_64 = _T_8156 % 5'h10; // @[util.scala 10:14:@4700.6]
  assign _T_8157 = _GEN_64[4:0]; // @[util.scala 10:14:@4700.6]
  assign _GEN_1120 = _T_8153 ? _T_8157 : {{1'd0}, head}; // @[StoreQueue.scala 229:50:@4698.4]
  assign _GEN_1234 = {{2'd0}, io_bbNumStores}; // @[util.scala 10:8:@4704.6]
  assign _T_8159 = tail + _GEN_1234; // @[util.scala 10:8:@4704.6]
  assign _GEN_65 = _T_8159 % 5'h10; // @[util.scala 10:14:@4705.6]
  assign _T_8160 = _GEN_65[4:0]; // @[util.scala 10:14:@4705.6]
  assign _GEN_1121 = io_bbStart ? _T_8160 : {{1'd0}, tail}; // @[StoreQueue.scala 233:20:@4703.4]
  assign _T_8162 = allocatedEntries_0 == 1'h0; // @[StoreQueue.scala 237:84:@4708.4]
  assign _T_8163 = storeCompleted_0 | _T_8162; // @[StoreQueue.scala 237:81:@4709.4]
  assign _T_8165 = allocatedEntries_1 == 1'h0; // @[StoreQueue.scala 237:84:@4710.4]
  assign _T_8166 = storeCompleted_1 | _T_8165; // @[StoreQueue.scala 237:81:@4711.4]
  assign _T_8168 = allocatedEntries_2 == 1'h0; // @[StoreQueue.scala 237:84:@4712.4]
  assign _T_8169 = storeCompleted_2 | _T_8168; // @[StoreQueue.scala 237:81:@4713.4]
  assign _T_8171 = allocatedEntries_3 == 1'h0; // @[StoreQueue.scala 237:84:@4714.4]
  assign _T_8172 = storeCompleted_3 | _T_8171; // @[StoreQueue.scala 237:81:@4715.4]
  assign _T_8174 = allocatedEntries_4 == 1'h0; // @[StoreQueue.scala 237:84:@4716.4]
  assign _T_8175 = storeCompleted_4 | _T_8174; // @[StoreQueue.scala 237:81:@4717.4]
  assign _T_8177 = allocatedEntries_5 == 1'h0; // @[StoreQueue.scala 237:84:@4718.4]
  assign _T_8178 = storeCompleted_5 | _T_8177; // @[StoreQueue.scala 237:81:@4719.4]
  assign _T_8180 = allocatedEntries_6 == 1'h0; // @[StoreQueue.scala 237:84:@4720.4]
  assign _T_8181 = storeCompleted_6 | _T_8180; // @[StoreQueue.scala 237:81:@4721.4]
  assign _T_8183 = allocatedEntries_7 == 1'h0; // @[StoreQueue.scala 237:84:@4722.4]
  assign _T_8184 = storeCompleted_7 | _T_8183; // @[StoreQueue.scala 237:81:@4723.4]
  assign _T_8186 = allocatedEntries_8 == 1'h0; // @[StoreQueue.scala 237:84:@4724.4]
  assign _T_8187 = storeCompleted_8 | _T_8186; // @[StoreQueue.scala 237:81:@4725.4]
  assign _T_8189 = allocatedEntries_9 == 1'h0; // @[StoreQueue.scala 237:84:@4726.4]
  assign _T_8190 = storeCompleted_9 | _T_8189; // @[StoreQueue.scala 237:81:@4727.4]
  assign _T_8192 = allocatedEntries_10 == 1'h0; // @[StoreQueue.scala 237:84:@4728.4]
  assign _T_8193 = storeCompleted_10 | _T_8192; // @[StoreQueue.scala 237:81:@4729.4]
  assign _T_8195 = allocatedEntries_11 == 1'h0; // @[StoreQueue.scala 237:84:@4730.4]
  assign _T_8196 = storeCompleted_11 | _T_8195; // @[StoreQueue.scala 237:81:@4731.4]
  assign _T_8198 = allocatedEntries_12 == 1'h0; // @[StoreQueue.scala 237:84:@4732.4]
  assign _T_8199 = storeCompleted_12 | _T_8198; // @[StoreQueue.scala 237:81:@4733.4]
  assign _T_8201 = allocatedEntries_13 == 1'h0; // @[StoreQueue.scala 237:84:@4734.4]
  assign _T_8202 = storeCompleted_13 | _T_8201; // @[StoreQueue.scala 237:81:@4735.4]
  assign _T_8204 = allocatedEntries_14 == 1'h0; // @[StoreQueue.scala 237:84:@4736.4]
  assign _T_8205 = storeCompleted_14 | _T_8204; // @[StoreQueue.scala 237:81:@4737.4]
  assign _T_8207 = allocatedEntries_15 == 1'h0; // @[StoreQueue.scala 237:84:@4738.4]
  assign _T_8208 = storeCompleted_15 | _T_8207; // @[StoreQueue.scala 237:81:@4739.4]
  assign _T_8233 = _T_8163 & _T_8166; // @[StoreQueue.scala 237:98:@4758.4]
  assign _T_8234 = _T_8233 & _T_8169; // @[StoreQueue.scala 237:98:@4759.4]
  assign _T_8235 = _T_8234 & _T_8172; // @[StoreQueue.scala 237:98:@4760.4]
  assign _T_8236 = _T_8235 & _T_8175; // @[StoreQueue.scala 237:98:@4761.4]
  assign _T_8237 = _T_8236 & _T_8178; // @[StoreQueue.scala 237:98:@4762.4]
  assign _T_8238 = _T_8237 & _T_8181; // @[StoreQueue.scala 237:98:@4763.4]
  assign _T_8239 = _T_8238 & _T_8184; // @[StoreQueue.scala 237:98:@4764.4]
  assign _T_8240 = _T_8239 & _T_8187; // @[StoreQueue.scala 237:98:@4765.4]
  assign _T_8241 = _T_8240 & _T_8190; // @[StoreQueue.scala 237:98:@4766.4]
  assign _T_8242 = _T_8241 & _T_8193; // @[StoreQueue.scala 237:98:@4767.4]
  assign _T_8243 = _T_8242 & _T_8196; // @[StoreQueue.scala 237:98:@4768.4]
  assign _T_8244 = _T_8243 & _T_8199; // @[StoreQueue.scala 237:98:@4769.4]
  assign _T_8245 = _T_8244 & _T_8202; // @[StoreQueue.scala 237:98:@4770.4]
  assign _T_8246 = _T_8245 & _T_8205; // @[StoreQueue.scala 237:98:@4771.4]
  assign _GEN_1123 = 4'h1 == head ? dataQ_1 : dataQ_0; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1124 = 4'h2 == head ? dataQ_2 : _GEN_1123; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1125 = 4'h3 == head ? dataQ_3 : _GEN_1124; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1126 = 4'h4 == head ? dataQ_4 : _GEN_1125; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1127 = 4'h5 == head ? dataQ_5 : _GEN_1126; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1128 = 4'h6 == head ? dataQ_6 : _GEN_1127; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1129 = 4'h7 == head ? dataQ_7 : _GEN_1128; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1130 = 4'h8 == head ? dataQ_8 : _GEN_1129; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1131 = 4'h9 == head ? dataQ_9 : _GEN_1130; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1132 = 4'ha == head ? dataQ_10 : _GEN_1131; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1133 = 4'hb == head ? dataQ_11 : _GEN_1132; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1134 = 4'hc == head ? dataQ_12 : _GEN_1133; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1135 = 4'hd == head ? dataQ_13 : _GEN_1134; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1136 = 4'he == head ? dataQ_14 : _GEN_1135; // @[StoreQueue.scala 252:21:@4841.4]
  assign io_storeTail = tail; // @[StoreQueue.scala 246:16:@4775.4]
  assign io_storeHead = head; // @[StoreQueue.scala 245:16:@4774.4]
  assign io_storeEmpty = _T_8246 & _T_8208; // @[StoreQueue.scala 237:17:@4773.4]
  assign io_storeAddrDone_0 = addrKnown_0; // @[StoreQueue.scala 250:20:@4824.4]
  assign io_storeAddrDone_1 = addrKnown_1; // @[StoreQueue.scala 250:20:@4825.4]
  assign io_storeAddrDone_2 = addrKnown_2; // @[StoreQueue.scala 250:20:@4826.4]
  assign io_storeAddrDone_3 = addrKnown_3; // @[StoreQueue.scala 250:20:@4827.4]
  assign io_storeAddrDone_4 = addrKnown_4; // @[StoreQueue.scala 250:20:@4828.4]
  assign io_storeAddrDone_5 = addrKnown_5; // @[StoreQueue.scala 250:20:@4829.4]
  assign io_storeAddrDone_6 = addrKnown_6; // @[StoreQueue.scala 250:20:@4830.4]
  assign io_storeAddrDone_7 = addrKnown_7; // @[StoreQueue.scala 250:20:@4831.4]
  assign io_storeAddrDone_8 = addrKnown_8; // @[StoreQueue.scala 250:20:@4832.4]
  assign io_storeAddrDone_9 = addrKnown_9; // @[StoreQueue.scala 250:20:@4833.4]
  assign io_storeAddrDone_10 = addrKnown_10; // @[StoreQueue.scala 250:20:@4834.4]
  assign io_storeAddrDone_11 = addrKnown_11; // @[StoreQueue.scala 250:20:@4835.4]
  assign io_storeAddrDone_12 = addrKnown_12; // @[StoreQueue.scala 250:20:@4836.4]
  assign io_storeAddrDone_13 = addrKnown_13; // @[StoreQueue.scala 250:20:@4837.4]
  assign io_storeAddrDone_14 = addrKnown_14; // @[StoreQueue.scala 250:20:@4838.4]
  assign io_storeAddrDone_15 = addrKnown_15; // @[StoreQueue.scala 250:20:@4839.4]
  assign io_storeDataDone_0 = dataKnown_0; // @[StoreQueue.scala 249:20:@4808.4]
  assign io_storeDataDone_1 = dataKnown_1; // @[StoreQueue.scala 249:20:@4809.4]
  assign io_storeDataDone_2 = dataKnown_2; // @[StoreQueue.scala 249:20:@4810.4]
  assign io_storeDataDone_3 = dataKnown_3; // @[StoreQueue.scala 249:20:@4811.4]
  assign io_storeDataDone_4 = dataKnown_4; // @[StoreQueue.scala 249:20:@4812.4]
  assign io_storeDataDone_5 = dataKnown_5; // @[StoreQueue.scala 249:20:@4813.4]
  assign io_storeDataDone_6 = dataKnown_6; // @[StoreQueue.scala 249:20:@4814.4]
  assign io_storeDataDone_7 = dataKnown_7; // @[StoreQueue.scala 249:20:@4815.4]
  assign io_storeDataDone_8 = dataKnown_8; // @[StoreQueue.scala 249:20:@4816.4]
  assign io_storeDataDone_9 = dataKnown_9; // @[StoreQueue.scala 249:20:@4817.4]
  assign io_storeDataDone_10 = dataKnown_10; // @[StoreQueue.scala 249:20:@4818.4]
  assign io_storeDataDone_11 = dataKnown_11; // @[StoreQueue.scala 249:20:@4819.4]
  assign io_storeDataDone_12 = dataKnown_12; // @[StoreQueue.scala 249:20:@4820.4]
  assign io_storeDataDone_13 = dataKnown_13; // @[StoreQueue.scala 249:20:@4821.4]
  assign io_storeDataDone_14 = dataKnown_14; // @[StoreQueue.scala 249:20:@4822.4]
  assign io_storeDataDone_15 = dataKnown_15; // @[StoreQueue.scala 249:20:@4823.4]
  assign io_storeAddrQueue_0 = addrQ_0; // @[StoreQueue.scala 247:21:@4776.4]
  assign io_storeAddrQueue_1 = addrQ_1; // @[StoreQueue.scala 247:21:@4777.4]
  assign io_storeAddrQueue_2 = addrQ_2; // @[StoreQueue.scala 247:21:@4778.4]
  assign io_storeAddrQueue_3 = addrQ_3; // @[StoreQueue.scala 247:21:@4779.4]
  assign io_storeAddrQueue_4 = addrQ_4; // @[StoreQueue.scala 247:21:@4780.4]
  assign io_storeAddrQueue_5 = addrQ_5; // @[StoreQueue.scala 247:21:@4781.4]
  assign io_storeAddrQueue_6 = addrQ_6; // @[StoreQueue.scala 247:21:@4782.4]
  assign io_storeAddrQueue_7 = addrQ_7; // @[StoreQueue.scala 247:21:@4783.4]
  assign io_storeAddrQueue_8 = addrQ_8; // @[StoreQueue.scala 247:21:@4784.4]
  assign io_storeAddrQueue_9 = addrQ_9; // @[StoreQueue.scala 247:21:@4785.4]
  assign io_storeAddrQueue_10 = addrQ_10; // @[StoreQueue.scala 247:21:@4786.4]
  assign io_storeAddrQueue_11 = addrQ_11; // @[StoreQueue.scala 247:21:@4787.4]
  assign io_storeAddrQueue_12 = addrQ_12; // @[StoreQueue.scala 247:21:@4788.4]
  assign io_storeAddrQueue_13 = addrQ_13; // @[StoreQueue.scala 247:21:@4789.4]
  assign io_storeAddrQueue_14 = addrQ_14; // @[StoreQueue.scala 247:21:@4790.4]
  assign io_storeAddrQueue_15 = addrQ_15; // @[StoreQueue.scala 247:21:@4791.4]
  assign io_storeDataQueue_0 = dataQ_0; // @[StoreQueue.scala 248:21:@4792.4]
  assign io_storeDataQueue_1 = dataQ_1; // @[StoreQueue.scala 248:21:@4793.4]
  assign io_storeDataQueue_2 = dataQ_2; // @[StoreQueue.scala 248:21:@4794.4]
  assign io_storeDataQueue_3 = dataQ_3; // @[StoreQueue.scala 248:21:@4795.4]
  assign io_storeDataQueue_4 = dataQ_4; // @[StoreQueue.scala 248:21:@4796.4]
  assign io_storeDataQueue_5 = dataQ_5; // @[StoreQueue.scala 248:21:@4797.4]
  assign io_storeDataQueue_6 = dataQ_6; // @[StoreQueue.scala 248:21:@4798.4]
  assign io_storeDataQueue_7 = dataQ_7; // @[StoreQueue.scala 248:21:@4799.4]
  assign io_storeDataQueue_8 = dataQ_8; // @[StoreQueue.scala 248:21:@4800.4]
  assign io_storeDataQueue_9 = dataQ_9; // @[StoreQueue.scala 248:21:@4801.4]
  assign io_storeDataQueue_10 = dataQ_10; // @[StoreQueue.scala 248:21:@4802.4]
  assign io_storeDataQueue_11 = dataQ_11; // @[StoreQueue.scala 248:21:@4803.4]
  assign io_storeDataQueue_12 = dataQ_12; // @[StoreQueue.scala 248:21:@4804.4]
  assign io_storeDataQueue_13 = dataQ_13; // @[StoreQueue.scala 248:21:@4805.4]
  assign io_storeDataQueue_14 = dataQ_14; // @[StoreQueue.scala 248:21:@4806.4]
  assign io_storeDataQueue_15 = dataQ_15; // @[StoreQueue.scala 248:21:@4807.4]
  assign io_storeAddrToMem = 4'hf == head ? addrQ_15 : _GEN_910; // @[StoreQueue.scala 253:21:@4842.4]
  assign io_storeDataToMem = 4'hf == head ? dataQ_15 : _GEN_1136; // @[StoreQueue.scala 252:21:@4841.4]
  assign io_storeEnableToMem = _T_3525 & _T_3542; // @[StoreQueue.scala 251:23:@4840.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  offsetQ_0 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  offsetQ_1 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  offsetQ_2 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  offsetQ_3 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  offsetQ_4 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  offsetQ_5 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  offsetQ_6 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  offsetQ_7 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  offsetQ_8 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  offsetQ_9 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  offsetQ_10 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  offsetQ_11 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  offsetQ_12 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  offsetQ_13 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  offsetQ_14 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  offsetQ_15 = _RAND_17[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  portQ_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  portQ_1 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  portQ_2 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  portQ_3 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  portQ_4 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  portQ_5 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  portQ_6 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  portQ_7 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  portQ_8 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  portQ_9 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  portQ_10 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  portQ_11 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  portQ_12 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  portQ_13 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  portQ_14 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  portQ_15 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  addrQ_0 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  addrQ_1 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  addrQ_2 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  addrQ_3 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  addrQ_4 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  addrQ_5 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  addrQ_6 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  addrQ_7 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  addrQ_8 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  addrQ_9 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  addrQ_10 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  addrQ_11 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  addrQ_12 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  addrQ_13 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  addrQ_14 = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  addrQ_15 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  dataQ_0 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  dataQ_1 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  dataQ_2 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  dataQ_3 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  dataQ_4 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  dataQ_5 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  dataQ_6 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  dataQ_7 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  dataQ_8 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  dataQ_9 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  dataQ_10 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  dataQ_11 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  dataQ_12 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  dataQ_13 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  dataQ_14 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  dataQ_15 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  addrKnown_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  addrKnown_1 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  addrKnown_2 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  addrKnown_3 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  addrKnown_4 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  addrKnown_5 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  addrKnown_6 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  addrKnown_7 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  addrKnown_8 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  addrKnown_9 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  addrKnown_10 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  addrKnown_11 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  addrKnown_12 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  addrKnown_13 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  addrKnown_14 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  addrKnown_15 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  dataKnown_0 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  dataKnown_1 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  dataKnown_2 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  dataKnown_3 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  dataKnown_4 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  dataKnown_5 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  dataKnown_6 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  dataKnown_7 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  dataKnown_8 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  dataKnown_9 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  dataKnown_10 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  dataKnown_11 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  dataKnown_12 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  dataKnown_13 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  dataKnown_14 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  dataKnown_15 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  allocatedEntries_0 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  allocatedEntries_1 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  allocatedEntries_2 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  allocatedEntries_3 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  allocatedEntries_4 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  allocatedEntries_5 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  allocatedEntries_6 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  allocatedEntries_7 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  allocatedEntries_8 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  allocatedEntries_9 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  allocatedEntries_10 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  allocatedEntries_11 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  allocatedEntries_12 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  allocatedEntries_13 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  allocatedEntries_14 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  allocatedEntries_15 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  storeCompleted_0 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  storeCompleted_1 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  storeCompleted_2 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  storeCompleted_3 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  storeCompleted_4 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  storeCompleted_5 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  storeCompleted_6 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  storeCompleted_7 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  storeCompleted_8 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  storeCompleted_9 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  storeCompleted_10 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  storeCompleted_11 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  storeCompleted_12 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  storeCompleted_13 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  storeCompleted_14 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  storeCompleted_15 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  checkBits_0 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  checkBits_1 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  checkBits_2 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  checkBits_3 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  checkBits_4 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  checkBits_5 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  checkBits_6 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  checkBits_7 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  checkBits_8 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  checkBits_9 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  checkBits_10 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  checkBits_11 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  checkBits_12 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  checkBits_13 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  checkBits_14 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  checkBits_15 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  previousLoadHead = _RAND_146[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      head <= 4'h0;
    end else begin
      head <= _GEN_1120[3:0];
    end
    if (reset) begin
      tail <= 4'h0;
    end else begin
      tail <= _GEN_1121[3:0];
    end
    if (reset) begin
      offsetQ_0 <= 4'h0;
    end else begin
      if (initBits_0) begin
        if (4'hf == _T_1804) begin
          offsetQ_0 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1804) begin
            offsetQ_0 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1804) begin
              offsetQ_0 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1804) begin
                offsetQ_0 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1804) begin
                  offsetQ_0 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1804) begin
                    offsetQ_0 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1804) begin
                      offsetQ_0 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1804) begin
                        offsetQ_0 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1804) begin
                          offsetQ_0 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1804) begin
                            offsetQ_0 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1804) begin
                              offsetQ_0 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1804) begin
                                offsetQ_0 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1804) begin
                                  offsetQ_0 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1804) begin
                                    offsetQ_0 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1804) begin
                                      offsetQ_0 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_0 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_1 <= 4'h0;
    end else begin
      if (initBits_1) begin
        if (4'hf == _T_1822) begin
          offsetQ_1 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1822) begin
            offsetQ_1 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1822) begin
              offsetQ_1 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1822) begin
                offsetQ_1 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1822) begin
                  offsetQ_1 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1822) begin
                    offsetQ_1 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1822) begin
                      offsetQ_1 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1822) begin
                        offsetQ_1 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1822) begin
                          offsetQ_1 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1822) begin
                            offsetQ_1 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1822) begin
                              offsetQ_1 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1822) begin
                                offsetQ_1 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1822) begin
                                  offsetQ_1 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1822) begin
                                    offsetQ_1 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1822) begin
                                      offsetQ_1 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_1 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_2 <= 4'h0;
    end else begin
      if (initBits_2) begin
        if (4'hf == _T_1840) begin
          offsetQ_2 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1840) begin
            offsetQ_2 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1840) begin
              offsetQ_2 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1840) begin
                offsetQ_2 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1840) begin
                  offsetQ_2 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1840) begin
                    offsetQ_2 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1840) begin
                      offsetQ_2 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1840) begin
                        offsetQ_2 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1840) begin
                          offsetQ_2 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1840) begin
                            offsetQ_2 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1840) begin
                              offsetQ_2 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1840) begin
                                offsetQ_2 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1840) begin
                                  offsetQ_2 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1840) begin
                                    offsetQ_2 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1840) begin
                                      offsetQ_2 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_2 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_3 <= 4'h0;
    end else begin
      if (initBits_3) begin
        if (4'hf == _T_1858) begin
          offsetQ_3 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1858) begin
            offsetQ_3 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1858) begin
              offsetQ_3 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1858) begin
                offsetQ_3 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1858) begin
                  offsetQ_3 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1858) begin
                    offsetQ_3 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1858) begin
                      offsetQ_3 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1858) begin
                        offsetQ_3 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1858) begin
                          offsetQ_3 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1858) begin
                            offsetQ_3 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1858) begin
                              offsetQ_3 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1858) begin
                                offsetQ_3 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1858) begin
                                  offsetQ_3 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1858) begin
                                    offsetQ_3 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1858) begin
                                      offsetQ_3 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_3 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_4 <= 4'h0;
    end else begin
      if (initBits_4) begin
        if (4'hf == _T_1876) begin
          offsetQ_4 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1876) begin
            offsetQ_4 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1876) begin
              offsetQ_4 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1876) begin
                offsetQ_4 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1876) begin
                  offsetQ_4 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1876) begin
                    offsetQ_4 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1876) begin
                      offsetQ_4 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1876) begin
                        offsetQ_4 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1876) begin
                          offsetQ_4 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1876) begin
                            offsetQ_4 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1876) begin
                              offsetQ_4 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1876) begin
                                offsetQ_4 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1876) begin
                                  offsetQ_4 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1876) begin
                                    offsetQ_4 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1876) begin
                                      offsetQ_4 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_4 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_5 <= 4'h0;
    end else begin
      if (initBits_5) begin
        if (4'hf == _T_1894) begin
          offsetQ_5 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1894) begin
            offsetQ_5 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1894) begin
              offsetQ_5 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1894) begin
                offsetQ_5 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1894) begin
                  offsetQ_5 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1894) begin
                    offsetQ_5 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1894) begin
                      offsetQ_5 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1894) begin
                        offsetQ_5 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1894) begin
                          offsetQ_5 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1894) begin
                            offsetQ_5 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1894) begin
                              offsetQ_5 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1894) begin
                                offsetQ_5 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1894) begin
                                  offsetQ_5 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1894) begin
                                    offsetQ_5 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1894) begin
                                      offsetQ_5 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_5 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_6 <= 4'h0;
    end else begin
      if (initBits_6) begin
        if (4'hf == _T_1912) begin
          offsetQ_6 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1912) begin
            offsetQ_6 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1912) begin
              offsetQ_6 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1912) begin
                offsetQ_6 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1912) begin
                  offsetQ_6 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1912) begin
                    offsetQ_6 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1912) begin
                      offsetQ_6 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1912) begin
                        offsetQ_6 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1912) begin
                          offsetQ_6 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1912) begin
                            offsetQ_6 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1912) begin
                              offsetQ_6 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1912) begin
                                offsetQ_6 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1912) begin
                                  offsetQ_6 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1912) begin
                                    offsetQ_6 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1912) begin
                                      offsetQ_6 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_6 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_7 <= 4'h0;
    end else begin
      if (initBits_7) begin
        if (4'hf == _T_1930) begin
          offsetQ_7 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1930) begin
            offsetQ_7 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1930) begin
              offsetQ_7 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1930) begin
                offsetQ_7 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1930) begin
                  offsetQ_7 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1930) begin
                    offsetQ_7 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1930) begin
                      offsetQ_7 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1930) begin
                        offsetQ_7 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1930) begin
                          offsetQ_7 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1930) begin
                            offsetQ_7 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1930) begin
                              offsetQ_7 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1930) begin
                                offsetQ_7 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1930) begin
                                  offsetQ_7 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1930) begin
                                    offsetQ_7 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1930) begin
                                      offsetQ_7 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_7 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_8 <= 4'h0;
    end else begin
      if (initBits_8) begin
        if (4'hf == _T_1948) begin
          offsetQ_8 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1948) begin
            offsetQ_8 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1948) begin
              offsetQ_8 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1948) begin
                offsetQ_8 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1948) begin
                  offsetQ_8 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1948) begin
                    offsetQ_8 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1948) begin
                      offsetQ_8 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1948) begin
                        offsetQ_8 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1948) begin
                          offsetQ_8 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1948) begin
                            offsetQ_8 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1948) begin
                              offsetQ_8 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1948) begin
                                offsetQ_8 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1948) begin
                                  offsetQ_8 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1948) begin
                                    offsetQ_8 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1948) begin
                                      offsetQ_8 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_8 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_9 <= 4'h0;
    end else begin
      if (initBits_9) begin
        if (4'hf == _T_1966) begin
          offsetQ_9 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1966) begin
            offsetQ_9 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1966) begin
              offsetQ_9 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1966) begin
                offsetQ_9 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1966) begin
                  offsetQ_9 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1966) begin
                    offsetQ_9 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1966) begin
                      offsetQ_9 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1966) begin
                        offsetQ_9 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1966) begin
                          offsetQ_9 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1966) begin
                            offsetQ_9 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1966) begin
                              offsetQ_9 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1966) begin
                                offsetQ_9 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1966) begin
                                  offsetQ_9 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1966) begin
                                    offsetQ_9 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1966) begin
                                      offsetQ_9 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_9 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_10 <= 4'h0;
    end else begin
      if (initBits_10) begin
        if (4'hf == _T_1984) begin
          offsetQ_10 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1984) begin
            offsetQ_10 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1984) begin
              offsetQ_10 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1984) begin
                offsetQ_10 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1984) begin
                  offsetQ_10 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1984) begin
                    offsetQ_10 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1984) begin
                      offsetQ_10 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1984) begin
                        offsetQ_10 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1984) begin
                          offsetQ_10 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1984) begin
                            offsetQ_10 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1984) begin
                              offsetQ_10 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1984) begin
                                offsetQ_10 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1984) begin
                                  offsetQ_10 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1984) begin
                                    offsetQ_10 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1984) begin
                                      offsetQ_10 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_10 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_11 <= 4'h0;
    end else begin
      if (initBits_11) begin
        if (4'hf == _T_2002) begin
          offsetQ_11 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2002) begin
            offsetQ_11 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2002) begin
              offsetQ_11 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2002) begin
                offsetQ_11 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2002) begin
                  offsetQ_11 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2002) begin
                    offsetQ_11 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2002) begin
                      offsetQ_11 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2002) begin
                        offsetQ_11 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2002) begin
                          offsetQ_11 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2002) begin
                            offsetQ_11 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2002) begin
                              offsetQ_11 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2002) begin
                                offsetQ_11 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2002) begin
                                  offsetQ_11 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2002) begin
                                    offsetQ_11 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2002) begin
                                      offsetQ_11 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_11 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_12 <= 4'h0;
    end else begin
      if (initBits_12) begin
        if (4'hf == _T_2020) begin
          offsetQ_12 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2020) begin
            offsetQ_12 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2020) begin
              offsetQ_12 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2020) begin
                offsetQ_12 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2020) begin
                  offsetQ_12 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2020) begin
                    offsetQ_12 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2020) begin
                      offsetQ_12 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2020) begin
                        offsetQ_12 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2020) begin
                          offsetQ_12 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2020) begin
                            offsetQ_12 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2020) begin
                              offsetQ_12 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2020) begin
                                offsetQ_12 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2020) begin
                                  offsetQ_12 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2020) begin
                                    offsetQ_12 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2020) begin
                                      offsetQ_12 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_12 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_13 <= 4'h0;
    end else begin
      if (initBits_13) begin
        if (4'hf == _T_2038) begin
          offsetQ_13 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2038) begin
            offsetQ_13 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2038) begin
              offsetQ_13 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2038) begin
                offsetQ_13 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2038) begin
                  offsetQ_13 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2038) begin
                    offsetQ_13 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2038) begin
                      offsetQ_13 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2038) begin
                        offsetQ_13 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2038) begin
                          offsetQ_13 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2038) begin
                            offsetQ_13 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2038) begin
                              offsetQ_13 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2038) begin
                                offsetQ_13 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2038) begin
                                  offsetQ_13 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2038) begin
                                    offsetQ_13 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2038) begin
                                      offsetQ_13 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_13 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_14 <= 4'h0;
    end else begin
      if (initBits_14) begin
        if (4'hf == _T_2056) begin
          offsetQ_14 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2056) begin
            offsetQ_14 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2056) begin
              offsetQ_14 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2056) begin
                offsetQ_14 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2056) begin
                  offsetQ_14 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2056) begin
                    offsetQ_14 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2056) begin
                      offsetQ_14 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2056) begin
                        offsetQ_14 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2056) begin
                          offsetQ_14 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2056) begin
                            offsetQ_14 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2056) begin
                              offsetQ_14 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2056) begin
                                offsetQ_14 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2056) begin
                                  offsetQ_14 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2056) begin
                                    offsetQ_14 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2056) begin
                                      offsetQ_14 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_14 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_15 <= 4'h0;
    end else begin
      if (initBits_15) begin
        if (4'hf == _T_2074) begin
          offsetQ_15 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2074) begin
            offsetQ_15 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2074) begin
              offsetQ_15 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2074) begin
                offsetQ_15 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2074) begin
                  offsetQ_15 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2074) begin
                    offsetQ_15 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2074) begin
                      offsetQ_15 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2074) begin
                        offsetQ_15 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2074) begin
                          offsetQ_15 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2074) begin
                            offsetQ_15 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2074) begin
                              offsetQ_15 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2074) begin
                                offsetQ_15 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2074) begin
                                  offsetQ_15 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2074) begin
                                    offsetQ_15 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2074) begin
                                      offsetQ_15 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_15 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        portQ_0 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        portQ_1 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        portQ_2 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        portQ_3 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        portQ_4 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        portQ_5 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        portQ_6 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        portQ_7 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        portQ_8 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        portQ_9 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        portQ_10 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        portQ_11 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        portQ_12 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        portQ_13 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        portQ_14 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        portQ_15 <= 1'h0;
      end
    end
    if (reset) begin
      addrQ_0 <= 32'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_7582) begin
          addrQ_0 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_1 <= 32'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_7618) begin
          addrQ_1 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_2 <= 32'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_7654) begin
          addrQ_2 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_3 <= 32'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_7690) begin
          addrQ_3 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_4 <= 32'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_7726) begin
          addrQ_4 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_5 <= 32'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_7762) begin
          addrQ_5 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_6 <= 32'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_7798) begin
          addrQ_6 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_7 <= 32'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_7834) begin
          addrQ_7 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_8 <= 32'h0;
    end else begin
      if (!(initBits_8)) begin
        if (_T_7870) begin
          addrQ_8 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_9 <= 32'h0;
    end else begin
      if (!(initBits_9)) begin
        if (_T_7906) begin
          addrQ_9 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_10 <= 32'h0;
    end else begin
      if (!(initBits_10)) begin
        if (_T_7942) begin
          addrQ_10 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_11 <= 32'h0;
    end else begin
      if (!(initBits_11)) begin
        if (_T_7978) begin
          addrQ_11 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_12 <= 32'h0;
    end else begin
      if (!(initBits_12)) begin
        if (_T_8014) begin
          addrQ_12 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_13 <= 32'h0;
    end else begin
      if (!(initBits_13)) begin
        if (_T_8050) begin
          addrQ_13 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_14 <= 32'h0;
    end else begin
      if (!(initBits_14)) begin
        if (_T_8086) begin
          addrQ_14 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_15 <= 32'h0;
    end else begin
      if (!(initBits_15)) begin
        if (_T_8122) begin
          addrQ_15 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_0 <= 32'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_7599) begin
          dataQ_0 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_1 <= 32'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_7635) begin
          dataQ_1 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_2 <= 32'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_7671) begin
          dataQ_2 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_3 <= 32'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_7707) begin
          dataQ_3 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_4 <= 32'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_7743) begin
          dataQ_4 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_5 <= 32'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_7779) begin
          dataQ_5 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_6 <= 32'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_7815) begin
          dataQ_6 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_7 <= 32'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_7851) begin
          dataQ_7 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_8 <= 32'h0;
    end else begin
      if (!(initBits_8)) begin
        if (_T_7887) begin
          dataQ_8 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_9 <= 32'h0;
    end else begin
      if (!(initBits_9)) begin
        if (_T_7923) begin
          dataQ_9 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_10 <= 32'h0;
    end else begin
      if (!(initBits_10)) begin
        if (_T_7959) begin
          dataQ_10 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_11 <= 32'h0;
    end else begin
      if (!(initBits_11)) begin
        if (_T_7995) begin
          dataQ_11 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_12 <= 32'h0;
    end else begin
      if (!(initBits_12)) begin
        if (_T_8031) begin
          dataQ_12 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_13 <= 32'h0;
    end else begin
      if (!(initBits_13)) begin
        if (_T_8067) begin
          dataQ_13 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_14 <= 32'h0;
    end else begin
      if (!(initBits_14)) begin
        if (_T_8103) begin
          dataQ_14 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_15 <= 32'h0;
    end else begin
      if (!(initBits_15)) begin
        if (_T_8139) begin
          dataQ_15 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        addrKnown_0 <= 1'h0;
      end else begin
        if (_T_7582) begin
          addrKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        addrKnown_1 <= 1'h0;
      end else begin
        if (_T_7618) begin
          addrKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        addrKnown_2 <= 1'h0;
      end else begin
        if (_T_7654) begin
          addrKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        addrKnown_3 <= 1'h0;
      end else begin
        if (_T_7690) begin
          addrKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        addrKnown_4 <= 1'h0;
      end else begin
        if (_T_7726) begin
          addrKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        addrKnown_5 <= 1'h0;
      end else begin
        if (_T_7762) begin
          addrKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        addrKnown_6 <= 1'h0;
      end else begin
        if (_T_7798) begin
          addrKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        addrKnown_7 <= 1'h0;
      end else begin
        if (_T_7834) begin
          addrKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        addrKnown_8 <= 1'h0;
      end else begin
        if (_T_7870) begin
          addrKnown_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        addrKnown_9 <= 1'h0;
      end else begin
        if (_T_7906) begin
          addrKnown_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        addrKnown_10 <= 1'h0;
      end else begin
        if (_T_7942) begin
          addrKnown_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        addrKnown_11 <= 1'h0;
      end else begin
        if (_T_7978) begin
          addrKnown_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        addrKnown_12 <= 1'h0;
      end else begin
        if (_T_8014) begin
          addrKnown_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        addrKnown_13 <= 1'h0;
      end else begin
        if (_T_8050) begin
          addrKnown_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        addrKnown_14 <= 1'h0;
      end else begin
        if (_T_8086) begin
          addrKnown_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        addrKnown_15 <= 1'h0;
      end else begin
        if (_T_8122) begin
          addrKnown_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        dataKnown_0 <= 1'h0;
      end else begin
        if (_T_7599) begin
          dataKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        dataKnown_1 <= 1'h0;
      end else begin
        if (_T_7635) begin
          dataKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        dataKnown_2 <= 1'h0;
      end else begin
        if (_T_7671) begin
          dataKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        dataKnown_3 <= 1'h0;
      end else begin
        if (_T_7707) begin
          dataKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        dataKnown_4 <= 1'h0;
      end else begin
        if (_T_7743) begin
          dataKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        dataKnown_5 <= 1'h0;
      end else begin
        if (_T_7779) begin
          dataKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        dataKnown_6 <= 1'h0;
      end else begin
        if (_T_7815) begin
          dataKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        dataKnown_7 <= 1'h0;
      end else begin
        if (_T_7851) begin
          dataKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        dataKnown_8 <= 1'h0;
      end else begin
        if (_T_7887) begin
          dataKnown_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        dataKnown_9 <= 1'h0;
      end else begin
        if (_T_7923) begin
          dataKnown_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        dataKnown_10 <= 1'h0;
      end else begin
        if (_T_7959) begin
          dataKnown_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        dataKnown_11 <= 1'h0;
      end else begin
        if (_T_7995) begin
          dataKnown_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        dataKnown_12 <= 1'h0;
      end else begin
        if (_T_8031) begin
          dataKnown_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        dataKnown_13 <= 1'h0;
      end else begin
        if (_T_8067) begin
          dataKnown_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        dataKnown_14 <= 1'h0;
      end else begin
        if (_T_8103) begin
          dataKnown_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        dataKnown_15 <= 1'h0;
      end else begin
        if (_T_8139) begin
          dataKnown_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      allocatedEntries_0 <= 1'h0;
    end else begin
      allocatedEntries_0 <= _T_1758;
    end
    if (reset) begin
      allocatedEntries_1 <= 1'h0;
    end else begin
      allocatedEntries_1 <= _T_1759;
    end
    if (reset) begin
      allocatedEntries_2 <= 1'h0;
    end else begin
      allocatedEntries_2 <= _T_1760;
    end
    if (reset) begin
      allocatedEntries_3 <= 1'h0;
    end else begin
      allocatedEntries_3 <= _T_1761;
    end
    if (reset) begin
      allocatedEntries_4 <= 1'h0;
    end else begin
      allocatedEntries_4 <= _T_1762;
    end
    if (reset) begin
      allocatedEntries_5 <= 1'h0;
    end else begin
      allocatedEntries_5 <= _T_1763;
    end
    if (reset) begin
      allocatedEntries_6 <= 1'h0;
    end else begin
      allocatedEntries_6 <= _T_1764;
    end
    if (reset) begin
      allocatedEntries_7 <= 1'h0;
    end else begin
      allocatedEntries_7 <= _T_1765;
    end
    if (reset) begin
      allocatedEntries_8 <= 1'h0;
    end else begin
      allocatedEntries_8 <= _T_1766;
    end
    if (reset) begin
      allocatedEntries_9 <= 1'h0;
    end else begin
      allocatedEntries_9 <= _T_1767;
    end
    if (reset) begin
      allocatedEntries_10 <= 1'h0;
    end else begin
      allocatedEntries_10 <= _T_1768;
    end
    if (reset) begin
      allocatedEntries_11 <= 1'h0;
    end else begin
      allocatedEntries_11 <= _T_1769;
    end
    if (reset) begin
      allocatedEntries_12 <= 1'h0;
    end else begin
      allocatedEntries_12 <= _T_1770;
    end
    if (reset) begin
      allocatedEntries_13 <= 1'h0;
    end else begin
      allocatedEntries_13 <= _T_1771;
    end
    if (reset) begin
      allocatedEntries_14 <= 1'h0;
    end else begin
      allocatedEntries_14 <= _T_1772;
    end
    if (reset) begin
      allocatedEntries_15 <= 1'h0;
    end else begin
      allocatedEntries_15 <= _T_1773;
    end
    if (reset) begin
      storeCompleted_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        storeCompleted_0 <= 1'h0;
      end else begin
        if (_T_3547) begin
          storeCompleted_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        storeCompleted_1 <= 1'h0;
      end else begin
        if (_T_3553) begin
          storeCompleted_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        storeCompleted_2 <= 1'h0;
      end else begin
        if (_T_3559) begin
          storeCompleted_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        storeCompleted_3 <= 1'h0;
      end else begin
        if (_T_3565) begin
          storeCompleted_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        storeCompleted_4 <= 1'h0;
      end else begin
        if (_T_3571) begin
          storeCompleted_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        storeCompleted_5 <= 1'h0;
      end else begin
        if (_T_3577) begin
          storeCompleted_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        storeCompleted_6 <= 1'h0;
      end else begin
        if (_T_3583) begin
          storeCompleted_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        storeCompleted_7 <= 1'h0;
      end else begin
        if (_T_3589) begin
          storeCompleted_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        storeCompleted_8 <= 1'h0;
      end else begin
        if (_T_3595) begin
          storeCompleted_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        storeCompleted_9 <= 1'h0;
      end else begin
        if (_T_3601) begin
          storeCompleted_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        storeCompleted_10 <= 1'h0;
      end else begin
        if (_T_3607) begin
          storeCompleted_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        storeCompleted_11 <= 1'h0;
      end else begin
        if (_T_3613) begin
          storeCompleted_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        storeCompleted_12 <= 1'h0;
      end else begin
        if (_T_3619) begin
          storeCompleted_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        storeCompleted_13 <= 1'h0;
      end else begin
        if (_T_3625) begin
          storeCompleted_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        storeCompleted_14 <= 1'h0;
      end else begin
        if (_T_3631) begin
          storeCompleted_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        storeCompleted_15 <= 1'h0;
      end else begin
        if (_T_3637) begin
          storeCompleted_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      checkBits_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        checkBits_0 <= _T_2101;
      end else begin
        if (io_loadEmpty) begin
          checkBits_0 <= 1'h0;
        end else begin
          if (_T_2105) begin
            checkBits_0 <= 1'h0;
          end else begin
            if (_T_2113) begin
              checkBits_0 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        checkBits_1 <= _T_2131;
      end else begin
        if (io_loadEmpty) begin
          checkBits_1 <= 1'h0;
        end else begin
          if (_T_2135) begin
            checkBits_1 <= 1'h0;
          end else begin
            if (_T_2143) begin
              checkBits_1 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        checkBits_2 <= _T_2161;
      end else begin
        if (io_loadEmpty) begin
          checkBits_2 <= 1'h0;
        end else begin
          if (_T_2165) begin
            checkBits_2 <= 1'h0;
          end else begin
            if (_T_2173) begin
              checkBits_2 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        checkBits_3 <= _T_2191;
      end else begin
        if (io_loadEmpty) begin
          checkBits_3 <= 1'h0;
        end else begin
          if (_T_2195) begin
            checkBits_3 <= 1'h0;
          end else begin
            if (_T_2203) begin
              checkBits_3 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        checkBits_4 <= _T_2221;
      end else begin
        if (io_loadEmpty) begin
          checkBits_4 <= 1'h0;
        end else begin
          if (_T_2225) begin
            checkBits_4 <= 1'h0;
          end else begin
            if (_T_2233) begin
              checkBits_4 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        checkBits_5 <= _T_2251;
      end else begin
        if (io_loadEmpty) begin
          checkBits_5 <= 1'h0;
        end else begin
          if (_T_2255) begin
            checkBits_5 <= 1'h0;
          end else begin
            if (_T_2263) begin
              checkBits_5 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        checkBits_6 <= _T_2281;
      end else begin
        if (io_loadEmpty) begin
          checkBits_6 <= 1'h0;
        end else begin
          if (_T_2285) begin
            checkBits_6 <= 1'h0;
          end else begin
            if (_T_2293) begin
              checkBits_6 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        checkBits_7 <= _T_2311;
      end else begin
        if (io_loadEmpty) begin
          checkBits_7 <= 1'h0;
        end else begin
          if (_T_2315) begin
            checkBits_7 <= 1'h0;
          end else begin
            if (_T_2323) begin
              checkBits_7 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        checkBits_8 <= _T_2341;
      end else begin
        if (io_loadEmpty) begin
          checkBits_8 <= 1'h0;
        end else begin
          if (_T_2345) begin
            checkBits_8 <= 1'h0;
          end else begin
            if (_T_2353) begin
              checkBits_8 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        checkBits_9 <= _T_2371;
      end else begin
        if (io_loadEmpty) begin
          checkBits_9 <= 1'h0;
        end else begin
          if (_T_2375) begin
            checkBits_9 <= 1'h0;
          end else begin
            if (_T_2383) begin
              checkBits_9 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        checkBits_10 <= _T_2401;
      end else begin
        if (io_loadEmpty) begin
          checkBits_10 <= 1'h0;
        end else begin
          if (_T_2405) begin
            checkBits_10 <= 1'h0;
          end else begin
            if (_T_2413) begin
              checkBits_10 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        checkBits_11 <= _T_2431;
      end else begin
        if (io_loadEmpty) begin
          checkBits_11 <= 1'h0;
        end else begin
          if (_T_2435) begin
            checkBits_11 <= 1'h0;
          end else begin
            if (_T_2443) begin
              checkBits_11 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        checkBits_12 <= _T_2461;
      end else begin
        if (io_loadEmpty) begin
          checkBits_12 <= 1'h0;
        end else begin
          if (_T_2465) begin
            checkBits_12 <= 1'h0;
          end else begin
            if (_T_2473) begin
              checkBits_12 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        checkBits_13 <= _T_2491;
      end else begin
        if (io_loadEmpty) begin
          checkBits_13 <= 1'h0;
        end else begin
          if (_T_2495) begin
            checkBits_13 <= 1'h0;
          end else begin
            if (_T_2503) begin
              checkBits_13 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        checkBits_14 <= _T_2521;
      end else begin
        if (io_loadEmpty) begin
          checkBits_14 <= 1'h0;
        end else begin
          if (_T_2525) begin
            checkBits_14 <= 1'h0;
          end else begin
            if (_T_2533) begin
              checkBits_14 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        checkBits_15 <= _T_2551;
      end else begin
        if (io_loadEmpty) begin
          checkBits_15 <= 1'h0;
        end else begin
          if (_T_2555) begin
            checkBits_15 <= 1'h0;
          end else begin
            if (_T_2563) begin
              checkBits_15 <= 1'h0;
            end
          end
        end
      end
    end
    previousLoadHead <= io_loadHead;
  end
endmodule
module LOAD_QUEUE_LSQ_data( // @[:@4844.2]
  input         clock, // @[:@4845.4]
  input         reset, // @[:@4846.4]
  input         io_bbStart, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_0, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_1, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_2, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_3, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_4, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_5, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_6, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_7, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_8, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_9, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_10, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_11, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_12, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_13, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_14, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_15, // @[:@4847.4]
  input         io_bbLoadPorts_1, // @[:@4847.4]
  input  [1:0]  io_bbNumLoads, // @[:@4847.4]
  output [3:0]  io_loadTail, // @[:@4847.4]
  output [3:0]  io_loadHead, // @[:@4847.4]
  output        io_loadEmpty, // @[:@4847.4]
  input  [3:0]  io_storeTail, // @[:@4847.4]
  input  [3:0]  io_storeHead, // @[:@4847.4]
  input         io_storeEmpty, // @[:@4847.4]
  input         io_storeAddrDone_0, // @[:@4847.4]
  input         io_storeAddrDone_1, // @[:@4847.4]
  input         io_storeAddrDone_2, // @[:@4847.4]
  input         io_storeAddrDone_3, // @[:@4847.4]
  input         io_storeAddrDone_4, // @[:@4847.4]
  input         io_storeAddrDone_5, // @[:@4847.4]
  input         io_storeAddrDone_6, // @[:@4847.4]
  input         io_storeAddrDone_7, // @[:@4847.4]
  input         io_storeAddrDone_8, // @[:@4847.4]
  input         io_storeAddrDone_9, // @[:@4847.4]
  input         io_storeAddrDone_10, // @[:@4847.4]
  input         io_storeAddrDone_11, // @[:@4847.4]
  input         io_storeAddrDone_12, // @[:@4847.4]
  input         io_storeAddrDone_13, // @[:@4847.4]
  input         io_storeAddrDone_14, // @[:@4847.4]
  input         io_storeAddrDone_15, // @[:@4847.4]
  input         io_storeDataDone_0, // @[:@4847.4]
  input         io_storeDataDone_1, // @[:@4847.4]
  input         io_storeDataDone_2, // @[:@4847.4]
  input         io_storeDataDone_3, // @[:@4847.4]
  input         io_storeDataDone_4, // @[:@4847.4]
  input         io_storeDataDone_5, // @[:@4847.4]
  input         io_storeDataDone_6, // @[:@4847.4]
  input         io_storeDataDone_7, // @[:@4847.4]
  input         io_storeDataDone_8, // @[:@4847.4]
  input         io_storeDataDone_9, // @[:@4847.4]
  input         io_storeDataDone_10, // @[:@4847.4]
  input         io_storeDataDone_11, // @[:@4847.4]
  input         io_storeDataDone_12, // @[:@4847.4]
  input         io_storeDataDone_13, // @[:@4847.4]
  input         io_storeDataDone_14, // @[:@4847.4]
  input         io_storeDataDone_15, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_0, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_1, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_2, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_3, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_4, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_5, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_6, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_7, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_8, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_9, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_10, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_11, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_12, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_13, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_14, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_15, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_0, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_1, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_2, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_3, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_4, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_5, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_6, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_7, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_8, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_9, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_10, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_11, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_12, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_13, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_14, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_15, // @[:@4847.4]
  output        io_loadAddrDone_0, // @[:@4847.4]
  output        io_loadAddrDone_1, // @[:@4847.4]
  output        io_loadAddrDone_2, // @[:@4847.4]
  output        io_loadAddrDone_3, // @[:@4847.4]
  output        io_loadAddrDone_4, // @[:@4847.4]
  output        io_loadAddrDone_5, // @[:@4847.4]
  output        io_loadAddrDone_6, // @[:@4847.4]
  output        io_loadAddrDone_7, // @[:@4847.4]
  output        io_loadAddrDone_8, // @[:@4847.4]
  output        io_loadAddrDone_9, // @[:@4847.4]
  output        io_loadAddrDone_10, // @[:@4847.4]
  output        io_loadAddrDone_11, // @[:@4847.4]
  output        io_loadAddrDone_12, // @[:@4847.4]
  output        io_loadAddrDone_13, // @[:@4847.4]
  output        io_loadAddrDone_14, // @[:@4847.4]
  output        io_loadAddrDone_15, // @[:@4847.4]
  output        io_loadDataDone_0, // @[:@4847.4]
  output        io_loadDataDone_1, // @[:@4847.4]
  output        io_loadDataDone_2, // @[:@4847.4]
  output        io_loadDataDone_3, // @[:@4847.4]
  output        io_loadDataDone_4, // @[:@4847.4]
  output        io_loadDataDone_5, // @[:@4847.4]
  output        io_loadDataDone_6, // @[:@4847.4]
  output        io_loadDataDone_7, // @[:@4847.4]
  output        io_loadDataDone_8, // @[:@4847.4]
  output        io_loadDataDone_9, // @[:@4847.4]
  output        io_loadDataDone_10, // @[:@4847.4]
  output        io_loadDataDone_11, // @[:@4847.4]
  output        io_loadDataDone_12, // @[:@4847.4]
  output        io_loadDataDone_13, // @[:@4847.4]
  output        io_loadDataDone_14, // @[:@4847.4]
  output        io_loadDataDone_15, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_0, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_1, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_2, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_3, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_4, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_5, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_6, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_7, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_8, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_9, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_10, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_11, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_12, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_13, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_14, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_15, // @[:@4847.4]
  input         io_loadAddrEnable_0, // @[:@4847.4]
  input         io_loadAddrEnable_1, // @[:@4847.4]
  input  [31:0] io_addrFromLoadPorts_0, // @[:@4847.4]
  input  [31:0] io_addrFromLoadPorts_1, // @[:@4847.4]
  input         io_loadPorts_0_ready, // @[:@4847.4]
  output        io_loadPorts_0_valid, // @[:@4847.4]
  output [31:0] io_loadPorts_0_bits, // @[:@4847.4]
  input         io_loadPorts_1_ready, // @[:@4847.4]
  output        io_loadPorts_1_valid, // @[:@4847.4]
  output [31:0] io_loadPorts_1_bits, // @[:@4847.4]
  input  [31:0] io_loadDataFromMem, // @[:@4847.4]
  output [31:0] io_loadAddrToMem, // @[:@4847.4]
  output        io_loadEnableToMem, // @[:@4847.4]
  input         io_memIsReadyForLoads // @[:@4847.4]
);
  reg [3:0] head; // @[LoadQueue.scala 50:21:@4849.4]
  reg [31:0] _RAND_0;
  reg [3:0] tail; // @[LoadQueue.scala 51:21:@4850.4]
  reg [31:0] _RAND_1;
  reg [3:0] offsetQ_0; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_2;
  reg [3:0] offsetQ_1; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_3;
  reg [3:0] offsetQ_2; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_4;
  reg [3:0] offsetQ_3; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_5;
  reg [3:0] offsetQ_4; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_6;
  reg [3:0] offsetQ_5; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_7;
  reg [3:0] offsetQ_6; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_8;
  reg [3:0] offsetQ_7; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_9;
  reg [3:0] offsetQ_8; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_10;
  reg [3:0] offsetQ_9; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_11;
  reg [3:0] offsetQ_10; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_12;
  reg [3:0] offsetQ_11; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_13;
  reg [3:0] offsetQ_12; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_14;
  reg [3:0] offsetQ_13; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_15;
  reg [3:0] offsetQ_14; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_16;
  reg [3:0] offsetQ_15; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_17;
  reg  portQ_0; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_18;
  reg  portQ_1; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_19;
  reg  portQ_2; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_20;
  reg  portQ_3; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_21;
  reg  portQ_4; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_22;
  reg  portQ_5; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_23;
  reg  portQ_6; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_24;
  reg  portQ_7; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_25;
  reg  portQ_8; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_26;
  reg  portQ_9; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_27;
  reg  portQ_10; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_28;
  reg  portQ_11; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_29;
  reg  portQ_12; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_30;
  reg  portQ_13; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_31;
  reg  portQ_14; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_32;
  reg  portQ_15; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_33;
  reg [31:0] addrQ_0; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_34;
  reg [31:0] addrQ_1; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_35;
  reg [31:0] addrQ_2; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_36;
  reg [31:0] addrQ_3; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_37;
  reg [31:0] addrQ_4; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_38;
  reg [31:0] addrQ_5; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_39;
  reg [31:0] addrQ_6; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_40;
  reg [31:0] addrQ_7; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_41;
  reg [31:0] addrQ_8; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_42;
  reg [31:0] addrQ_9; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_43;
  reg [31:0] addrQ_10; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_44;
  reg [31:0] addrQ_11; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_45;
  reg [31:0] addrQ_12; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_46;
  reg [31:0] addrQ_13; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_47;
  reg [31:0] addrQ_14; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_48;
  reg [31:0] addrQ_15; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_49;
  reg [31:0] dataQ_0; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_50;
  reg [31:0] dataQ_1; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_51;
  reg [31:0] dataQ_2; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_52;
  reg [31:0] dataQ_3; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_53;
  reg [31:0] dataQ_4; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_54;
  reg [31:0] dataQ_5; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_55;
  reg [31:0] dataQ_6; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_56;
  reg [31:0] dataQ_7; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_57;
  reg [31:0] dataQ_8; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_58;
  reg [31:0] dataQ_9; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_59;
  reg [31:0] dataQ_10; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_60;
  reg [31:0] dataQ_11; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_61;
  reg [31:0] dataQ_12; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_62;
  reg [31:0] dataQ_13; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_63;
  reg [31:0] dataQ_14; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_64;
  reg [31:0] dataQ_15; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_65;
  reg  addrKnown_0; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_66;
  reg  addrKnown_1; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_67;
  reg  addrKnown_2; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_68;
  reg  addrKnown_3; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_69;
  reg  addrKnown_4; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_70;
  reg  addrKnown_5; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_71;
  reg  addrKnown_6; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_72;
  reg  addrKnown_7; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_73;
  reg  addrKnown_8; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_74;
  reg  addrKnown_9; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_75;
  reg  addrKnown_10; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_76;
  reg  addrKnown_11; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_77;
  reg  addrKnown_12; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_78;
  reg  addrKnown_13; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_79;
  reg  addrKnown_14; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_80;
  reg  addrKnown_15; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_81;
  reg  dataKnown_0; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_82;
  reg  dataKnown_1; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_83;
  reg  dataKnown_2; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_84;
  reg  dataKnown_3; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_85;
  reg  dataKnown_4; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_86;
  reg  dataKnown_5; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_87;
  reg  dataKnown_6; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_88;
  reg  dataKnown_7; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_89;
  reg  dataKnown_8; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_90;
  reg  dataKnown_9; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_91;
  reg  dataKnown_10; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_92;
  reg  dataKnown_11; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_93;
  reg  dataKnown_12; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_94;
  reg  dataKnown_13; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_95;
  reg  dataKnown_14; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_96;
  reg  dataKnown_15; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_97;
  reg  loadCompleted_0; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_98;
  reg  loadCompleted_1; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_99;
  reg  loadCompleted_2; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_100;
  reg  loadCompleted_3; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_101;
  reg  loadCompleted_4; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_102;
  reg  loadCompleted_5; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_103;
  reg  loadCompleted_6; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_104;
  reg  loadCompleted_7; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_105;
  reg  loadCompleted_8; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_106;
  reg  loadCompleted_9; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_107;
  reg  loadCompleted_10; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_108;
  reg  loadCompleted_11; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_109;
  reg  loadCompleted_12; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_110;
  reg  loadCompleted_13; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_111;
  reg  loadCompleted_14; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_112;
  reg  loadCompleted_15; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_113;
  reg  allocatedEntries_0; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_114;
  reg  allocatedEntries_1; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_115;
  reg  allocatedEntries_2; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_116;
  reg  allocatedEntries_3; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_117;
  reg  allocatedEntries_4; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_118;
  reg  allocatedEntries_5; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_119;
  reg  allocatedEntries_6; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_120;
  reg  allocatedEntries_7; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_121;
  reg  allocatedEntries_8; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_122;
  reg  allocatedEntries_9; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_123;
  reg  allocatedEntries_10; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_124;
  reg  allocatedEntries_11; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_125;
  reg  allocatedEntries_12; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_126;
  reg  allocatedEntries_13; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_127;
  reg  allocatedEntries_14; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_128;
  reg  allocatedEntries_15; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_129;
  reg  bypassInitiated_0; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_130;
  reg  bypassInitiated_1; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_131;
  reg  bypassInitiated_2; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_132;
  reg  bypassInitiated_3; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_133;
  reg  bypassInitiated_4; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_134;
  reg  bypassInitiated_5; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_135;
  reg  bypassInitiated_6; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_136;
  reg  bypassInitiated_7; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_137;
  reg  bypassInitiated_8; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_138;
  reg  bypassInitiated_9; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_139;
  reg  bypassInitiated_10; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_140;
  reg  bypassInitiated_11; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_141;
  reg  bypassInitiated_12; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_142;
  reg  bypassInitiated_13; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_143;
  reg  bypassInitiated_14; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_144;
  reg  bypassInitiated_15; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_145;
  reg  checkBits_0; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_146;
  reg  checkBits_1; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_147;
  reg  checkBits_2; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_148;
  reg  checkBits_3; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_149;
  reg  checkBits_4; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_150;
  reg  checkBits_5; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_151;
  reg  checkBits_6; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_152;
  reg  checkBits_7; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_153;
  reg  checkBits_8; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_154;
  reg  checkBits_9; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_155;
  reg  checkBits_10; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_156;
  reg  checkBits_11; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_157;
  reg  checkBits_12; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_158;
  reg  checkBits_13; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_159;
  reg  checkBits_14; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_160;
  reg  checkBits_15; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_161;
  wire [5:0] _GEN_2312; // @[util.scala 14:20:@5032.4]
  wire [6:0] _T_1724; // @[util.scala 14:20:@5032.4]
  wire [6:0] _T_1725; // @[util.scala 14:20:@5033.4]
  wire [5:0] _T_1726; // @[util.scala 14:20:@5034.4]
  wire [5:0] _GEN_0; // @[util.scala 14:25:@5035.4]
  wire [4:0] _T_1727; // @[util.scala 14:25:@5035.4]
  wire [4:0] _GEN_2313; // @[LoadQueue.scala 71:46:@5036.4]
  wire  _T_1728; // @[LoadQueue.scala 71:46:@5036.4]
  wire  initBits_0; // @[LoadQueue.scala 71:63:@5037.4]
  wire [6:0] _T_1733; // @[util.scala 14:20:@5039.4]
  wire [6:0] _T_1734; // @[util.scala 14:20:@5040.4]
  wire [5:0] _T_1735; // @[util.scala 14:20:@5041.4]
  wire [5:0] _GEN_16; // @[util.scala 14:25:@5042.4]
  wire [4:0] _T_1736; // @[util.scala 14:25:@5042.4]
  wire  _T_1737; // @[LoadQueue.scala 71:46:@5043.4]
  wire  initBits_1; // @[LoadQueue.scala 71:63:@5044.4]
  wire [6:0] _T_1742; // @[util.scala 14:20:@5046.4]
  wire [6:0] _T_1743; // @[util.scala 14:20:@5047.4]
  wire [5:0] _T_1744; // @[util.scala 14:20:@5048.4]
  wire [5:0] _GEN_34; // @[util.scala 14:25:@5049.4]
  wire [4:0] _T_1745; // @[util.scala 14:25:@5049.4]
  wire  _T_1746; // @[LoadQueue.scala 71:46:@5050.4]
  wire  initBits_2; // @[LoadQueue.scala 71:63:@5051.4]
  wire [6:0] _T_1751; // @[util.scala 14:20:@5053.4]
  wire [6:0] _T_1752; // @[util.scala 14:20:@5054.4]
  wire [5:0] _T_1753; // @[util.scala 14:20:@5055.4]
  wire [5:0] _GEN_50; // @[util.scala 14:25:@5056.4]
  wire [4:0] _T_1754; // @[util.scala 14:25:@5056.4]
  wire  _T_1755; // @[LoadQueue.scala 71:46:@5057.4]
  wire  initBits_3; // @[LoadQueue.scala 71:63:@5058.4]
  wire [6:0] _T_1760; // @[util.scala 14:20:@5060.4]
  wire [6:0] _T_1761; // @[util.scala 14:20:@5061.4]
  wire [5:0] _T_1762; // @[util.scala 14:20:@5062.4]
  wire [5:0] _GEN_68; // @[util.scala 14:25:@5063.4]
  wire [4:0] _T_1763; // @[util.scala 14:25:@5063.4]
  wire  _T_1764; // @[LoadQueue.scala 71:46:@5064.4]
  wire  initBits_4; // @[LoadQueue.scala 71:63:@5065.4]
  wire [6:0] _T_1769; // @[util.scala 14:20:@5067.4]
  wire [6:0] _T_1770; // @[util.scala 14:20:@5068.4]
  wire [5:0] _T_1771; // @[util.scala 14:20:@5069.4]
  wire [5:0] _GEN_84; // @[util.scala 14:25:@5070.4]
  wire [4:0] _T_1772; // @[util.scala 14:25:@5070.4]
  wire  _T_1773; // @[LoadQueue.scala 71:46:@5071.4]
  wire  initBits_5; // @[LoadQueue.scala 71:63:@5072.4]
  wire [6:0] _T_1778; // @[util.scala 14:20:@5074.4]
  wire [6:0] _T_1779; // @[util.scala 14:20:@5075.4]
  wire [5:0] _T_1780; // @[util.scala 14:20:@5076.4]
  wire [5:0] _GEN_102; // @[util.scala 14:25:@5077.4]
  wire [4:0] _T_1781; // @[util.scala 14:25:@5077.4]
  wire  _T_1782; // @[LoadQueue.scala 71:46:@5078.4]
  wire  initBits_6; // @[LoadQueue.scala 71:63:@5079.4]
  wire [6:0] _T_1787; // @[util.scala 14:20:@5081.4]
  wire [6:0] _T_1788; // @[util.scala 14:20:@5082.4]
  wire [5:0] _T_1789; // @[util.scala 14:20:@5083.4]
  wire [5:0] _GEN_118; // @[util.scala 14:25:@5084.4]
  wire [4:0] _T_1790; // @[util.scala 14:25:@5084.4]
  wire  _T_1791; // @[LoadQueue.scala 71:46:@5085.4]
  wire  initBits_7; // @[LoadQueue.scala 71:63:@5086.4]
  wire [6:0] _T_1796; // @[util.scala 14:20:@5088.4]
  wire [6:0] _T_1797; // @[util.scala 14:20:@5089.4]
  wire [5:0] _T_1798; // @[util.scala 14:20:@5090.4]
  wire [5:0] _GEN_136; // @[util.scala 14:25:@5091.4]
  wire [4:0] _T_1799; // @[util.scala 14:25:@5091.4]
  wire  _T_1800; // @[LoadQueue.scala 71:46:@5092.4]
  wire  initBits_8; // @[LoadQueue.scala 71:63:@5093.4]
  wire [6:0] _T_1805; // @[util.scala 14:20:@5095.4]
  wire [6:0] _T_1806; // @[util.scala 14:20:@5096.4]
  wire [5:0] _T_1807; // @[util.scala 14:20:@5097.4]
  wire [5:0] _GEN_152; // @[util.scala 14:25:@5098.4]
  wire [4:0] _T_1808; // @[util.scala 14:25:@5098.4]
  wire  _T_1809; // @[LoadQueue.scala 71:46:@5099.4]
  wire  initBits_9; // @[LoadQueue.scala 71:63:@5100.4]
  wire [6:0] _T_1814; // @[util.scala 14:20:@5102.4]
  wire [6:0] _T_1815; // @[util.scala 14:20:@5103.4]
  wire [5:0] _T_1816; // @[util.scala 14:20:@5104.4]
  wire [5:0] _GEN_170; // @[util.scala 14:25:@5105.4]
  wire [4:0] _T_1817; // @[util.scala 14:25:@5105.4]
  wire  _T_1818; // @[LoadQueue.scala 71:46:@5106.4]
  wire  initBits_10; // @[LoadQueue.scala 71:63:@5107.4]
  wire [6:0] _T_1823; // @[util.scala 14:20:@5109.4]
  wire [6:0] _T_1824; // @[util.scala 14:20:@5110.4]
  wire [5:0] _T_1825; // @[util.scala 14:20:@5111.4]
  wire [5:0] _GEN_186; // @[util.scala 14:25:@5112.4]
  wire [4:0] _T_1826; // @[util.scala 14:25:@5112.4]
  wire  _T_1827; // @[LoadQueue.scala 71:46:@5113.4]
  wire  initBits_11; // @[LoadQueue.scala 71:63:@5114.4]
  wire [6:0] _T_1832; // @[util.scala 14:20:@5116.4]
  wire [6:0] _T_1833; // @[util.scala 14:20:@5117.4]
  wire [5:0] _T_1834; // @[util.scala 14:20:@5118.4]
  wire [5:0] _GEN_204; // @[util.scala 14:25:@5119.4]
  wire [4:0] _T_1835; // @[util.scala 14:25:@5119.4]
  wire  _T_1836; // @[LoadQueue.scala 71:46:@5120.4]
  wire  initBits_12; // @[LoadQueue.scala 71:63:@5121.4]
  wire [6:0] _T_1841; // @[util.scala 14:20:@5123.4]
  wire [6:0] _T_1842; // @[util.scala 14:20:@5124.4]
  wire [5:0] _T_1843; // @[util.scala 14:20:@5125.4]
  wire [5:0] _GEN_220; // @[util.scala 14:25:@5126.4]
  wire [4:0] _T_1844; // @[util.scala 14:25:@5126.4]
  wire  _T_1845; // @[LoadQueue.scala 71:46:@5127.4]
  wire  initBits_13; // @[LoadQueue.scala 71:63:@5128.4]
  wire [6:0] _T_1850; // @[util.scala 14:20:@5130.4]
  wire [6:0] _T_1851; // @[util.scala 14:20:@5131.4]
  wire [5:0] _T_1852; // @[util.scala 14:20:@5132.4]
  wire [5:0] _GEN_238; // @[util.scala 14:25:@5133.4]
  wire [4:0] _T_1853; // @[util.scala 14:25:@5133.4]
  wire  _T_1854; // @[LoadQueue.scala 71:46:@5134.4]
  wire  initBits_14; // @[LoadQueue.scala 71:63:@5135.4]
  wire [6:0] _T_1859; // @[util.scala 14:20:@5137.4]
  wire [6:0] _T_1860; // @[util.scala 14:20:@5138.4]
  wire [5:0] _T_1861; // @[util.scala 14:20:@5139.4]
  wire [5:0] _GEN_254; // @[util.scala 14:25:@5140.4]
  wire [4:0] _T_1862; // @[util.scala 14:25:@5140.4]
  wire  _T_1863; // @[LoadQueue.scala 71:46:@5141.4]
  wire  initBits_15; // @[LoadQueue.scala 71:63:@5142.4]
  wire  _T_1886; // @[LoadQueue.scala 73:78:@5160.4]
  wire  _T_1887; // @[LoadQueue.scala 73:78:@5161.4]
  wire  _T_1888; // @[LoadQueue.scala 73:78:@5162.4]
  wire  _T_1889; // @[LoadQueue.scala 73:78:@5163.4]
  wire  _T_1890; // @[LoadQueue.scala 73:78:@5164.4]
  wire  _T_1891; // @[LoadQueue.scala 73:78:@5165.4]
  wire  _T_1892; // @[LoadQueue.scala 73:78:@5166.4]
  wire  _T_1893; // @[LoadQueue.scala 73:78:@5167.4]
  wire  _T_1894; // @[LoadQueue.scala 73:78:@5168.4]
  wire  _T_1895; // @[LoadQueue.scala 73:78:@5169.4]
  wire  _T_1896; // @[LoadQueue.scala 73:78:@5170.4]
  wire  _T_1897; // @[LoadQueue.scala 73:78:@5171.4]
  wire  _T_1898; // @[LoadQueue.scala 73:78:@5172.4]
  wire  _T_1899; // @[LoadQueue.scala 73:78:@5173.4]
  wire  _T_1900; // @[LoadQueue.scala 73:78:@5174.4]
  wire  _T_1901; // @[LoadQueue.scala 73:78:@5175.4]
  wire [3:0] _T_1932; // @[:@5215.6]
  wire [3:0] _GEN_1; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_2; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_3; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_4; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_5; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_6; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_7; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_8; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_9; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_10; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_11; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_12; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_13; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_14; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_15; // @[LoadQueue.scala 77:20:@5216.6]
  wire  _GEN_17; // @[LoadQueue.scala 78:18:@5223.6]
  wire  _GEN_18; // @[LoadQueue.scala 78:18:@5223.6]
  wire  _GEN_19; // @[LoadQueue.scala 78:18:@5223.6]
  wire  _GEN_20; // @[LoadQueue.scala 78:18:@5223.6]
  wire  _GEN_21; // @[LoadQueue.scala 78:18:@5223.6]
  wire  _GEN_22; // @[LoadQueue.scala 78:18:@5223.6]
  wire  _GEN_23; // @[LoadQueue.scala 78:18:@5223.6]
  wire  _GEN_24; // @[LoadQueue.scala 78:18:@5223.6]
  wire  _GEN_25; // @[LoadQueue.scala 78:18:@5223.6]
  wire  _GEN_26; // @[LoadQueue.scala 78:18:@5223.6]
  wire  _GEN_27; // @[LoadQueue.scala 78:18:@5223.6]
  wire  _GEN_28; // @[LoadQueue.scala 78:18:@5223.6]
  wire  _GEN_29; // @[LoadQueue.scala 78:18:@5223.6]
  wire  _GEN_30; // @[LoadQueue.scala 78:18:@5223.6]
  wire  _GEN_31; // @[LoadQueue.scala 78:18:@5223.6]
  wire [3:0] _GEN_32; // @[LoadQueue.scala 76:25:@5209.4]
  wire  _GEN_33; // @[LoadQueue.scala 76:25:@5209.4]
  wire [3:0] _T_1950; // @[:@5231.6]
  wire [3:0] _GEN_35; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_36; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_37; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_38; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_39; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_40; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_41; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_42; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_43; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_44; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_45; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_46; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_47; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_48; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_49; // @[LoadQueue.scala 77:20:@5232.6]
  wire  _GEN_51; // @[LoadQueue.scala 78:18:@5239.6]
  wire  _GEN_52; // @[LoadQueue.scala 78:18:@5239.6]
  wire  _GEN_53; // @[LoadQueue.scala 78:18:@5239.6]
  wire  _GEN_54; // @[LoadQueue.scala 78:18:@5239.6]
  wire  _GEN_55; // @[LoadQueue.scala 78:18:@5239.6]
  wire  _GEN_56; // @[LoadQueue.scala 78:18:@5239.6]
  wire  _GEN_57; // @[LoadQueue.scala 78:18:@5239.6]
  wire  _GEN_58; // @[LoadQueue.scala 78:18:@5239.6]
  wire  _GEN_59; // @[LoadQueue.scala 78:18:@5239.6]
  wire  _GEN_60; // @[LoadQueue.scala 78:18:@5239.6]
  wire  _GEN_61; // @[LoadQueue.scala 78:18:@5239.6]
  wire  _GEN_62; // @[LoadQueue.scala 78:18:@5239.6]
  wire  _GEN_63; // @[LoadQueue.scala 78:18:@5239.6]
  wire  _GEN_64; // @[LoadQueue.scala 78:18:@5239.6]
  wire  _GEN_65; // @[LoadQueue.scala 78:18:@5239.6]
  wire [3:0] _GEN_66; // @[LoadQueue.scala 76:25:@5225.4]
  wire  _GEN_67; // @[LoadQueue.scala 76:25:@5225.4]
  wire [3:0] _T_1968; // @[:@5247.6]
  wire [3:0] _GEN_69; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_70; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_71; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_72; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_73; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_74; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_75; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_76; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_77; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_78; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_79; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_80; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_81; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_82; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_83; // @[LoadQueue.scala 77:20:@5248.6]
  wire  _GEN_85; // @[LoadQueue.scala 78:18:@5255.6]
  wire  _GEN_86; // @[LoadQueue.scala 78:18:@5255.6]
  wire  _GEN_87; // @[LoadQueue.scala 78:18:@5255.6]
  wire  _GEN_88; // @[LoadQueue.scala 78:18:@5255.6]
  wire  _GEN_89; // @[LoadQueue.scala 78:18:@5255.6]
  wire  _GEN_90; // @[LoadQueue.scala 78:18:@5255.6]
  wire  _GEN_91; // @[LoadQueue.scala 78:18:@5255.6]
  wire  _GEN_92; // @[LoadQueue.scala 78:18:@5255.6]
  wire  _GEN_93; // @[LoadQueue.scala 78:18:@5255.6]
  wire  _GEN_94; // @[LoadQueue.scala 78:18:@5255.6]
  wire  _GEN_95; // @[LoadQueue.scala 78:18:@5255.6]
  wire  _GEN_96; // @[LoadQueue.scala 78:18:@5255.6]
  wire  _GEN_97; // @[LoadQueue.scala 78:18:@5255.6]
  wire  _GEN_98; // @[LoadQueue.scala 78:18:@5255.6]
  wire  _GEN_99; // @[LoadQueue.scala 78:18:@5255.6]
  wire [3:0] _GEN_100; // @[LoadQueue.scala 76:25:@5241.4]
  wire  _GEN_101; // @[LoadQueue.scala 76:25:@5241.4]
  wire [3:0] _T_1986; // @[:@5263.6]
  wire [3:0] _GEN_103; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_104; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_105; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_106; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_107; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_108; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_109; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_110; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_111; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_112; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_113; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_114; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_115; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_116; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_117; // @[LoadQueue.scala 77:20:@5264.6]
  wire  _GEN_119; // @[LoadQueue.scala 78:18:@5271.6]
  wire  _GEN_120; // @[LoadQueue.scala 78:18:@5271.6]
  wire  _GEN_121; // @[LoadQueue.scala 78:18:@5271.6]
  wire  _GEN_122; // @[LoadQueue.scala 78:18:@5271.6]
  wire  _GEN_123; // @[LoadQueue.scala 78:18:@5271.6]
  wire  _GEN_124; // @[LoadQueue.scala 78:18:@5271.6]
  wire  _GEN_125; // @[LoadQueue.scala 78:18:@5271.6]
  wire  _GEN_126; // @[LoadQueue.scala 78:18:@5271.6]
  wire  _GEN_127; // @[LoadQueue.scala 78:18:@5271.6]
  wire  _GEN_128; // @[LoadQueue.scala 78:18:@5271.6]
  wire  _GEN_129; // @[LoadQueue.scala 78:18:@5271.6]
  wire  _GEN_130; // @[LoadQueue.scala 78:18:@5271.6]
  wire  _GEN_131; // @[LoadQueue.scala 78:18:@5271.6]
  wire  _GEN_132; // @[LoadQueue.scala 78:18:@5271.6]
  wire  _GEN_133; // @[LoadQueue.scala 78:18:@5271.6]
  wire [3:0] _GEN_134; // @[LoadQueue.scala 76:25:@5257.4]
  wire  _GEN_135; // @[LoadQueue.scala 76:25:@5257.4]
  wire [3:0] _T_2004; // @[:@5279.6]
  wire [3:0] _GEN_137; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_138; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_139; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_140; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_141; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_142; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_143; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_144; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_145; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_146; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_147; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_148; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_149; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_150; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_151; // @[LoadQueue.scala 77:20:@5280.6]
  wire  _GEN_153; // @[LoadQueue.scala 78:18:@5287.6]
  wire  _GEN_154; // @[LoadQueue.scala 78:18:@5287.6]
  wire  _GEN_155; // @[LoadQueue.scala 78:18:@5287.6]
  wire  _GEN_156; // @[LoadQueue.scala 78:18:@5287.6]
  wire  _GEN_157; // @[LoadQueue.scala 78:18:@5287.6]
  wire  _GEN_158; // @[LoadQueue.scala 78:18:@5287.6]
  wire  _GEN_159; // @[LoadQueue.scala 78:18:@5287.6]
  wire  _GEN_160; // @[LoadQueue.scala 78:18:@5287.6]
  wire  _GEN_161; // @[LoadQueue.scala 78:18:@5287.6]
  wire  _GEN_162; // @[LoadQueue.scala 78:18:@5287.6]
  wire  _GEN_163; // @[LoadQueue.scala 78:18:@5287.6]
  wire  _GEN_164; // @[LoadQueue.scala 78:18:@5287.6]
  wire  _GEN_165; // @[LoadQueue.scala 78:18:@5287.6]
  wire  _GEN_166; // @[LoadQueue.scala 78:18:@5287.6]
  wire  _GEN_167; // @[LoadQueue.scala 78:18:@5287.6]
  wire [3:0] _GEN_168; // @[LoadQueue.scala 76:25:@5273.4]
  wire  _GEN_169; // @[LoadQueue.scala 76:25:@5273.4]
  wire [3:0] _T_2022; // @[:@5295.6]
  wire [3:0] _GEN_171; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_172; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_173; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_174; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_175; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_176; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_177; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_178; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_179; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_180; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_181; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_182; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_183; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_184; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_185; // @[LoadQueue.scala 77:20:@5296.6]
  wire  _GEN_187; // @[LoadQueue.scala 78:18:@5303.6]
  wire  _GEN_188; // @[LoadQueue.scala 78:18:@5303.6]
  wire  _GEN_189; // @[LoadQueue.scala 78:18:@5303.6]
  wire  _GEN_190; // @[LoadQueue.scala 78:18:@5303.6]
  wire  _GEN_191; // @[LoadQueue.scala 78:18:@5303.6]
  wire  _GEN_192; // @[LoadQueue.scala 78:18:@5303.6]
  wire  _GEN_193; // @[LoadQueue.scala 78:18:@5303.6]
  wire  _GEN_194; // @[LoadQueue.scala 78:18:@5303.6]
  wire  _GEN_195; // @[LoadQueue.scala 78:18:@5303.6]
  wire  _GEN_196; // @[LoadQueue.scala 78:18:@5303.6]
  wire  _GEN_197; // @[LoadQueue.scala 78:18:@5303.6]
  wire  _GEN_198; // @[LoadQueue.scala 78:18:@5303.6]
  wire  _GEN_199; // @[LoadQueue.scala 78:18:@5303.6]
  wire  _GEN_200; // @[LoadQueue.scala 78:18:@5303.6]
  wire  _GEN_201; // @[LoadQueue.scala 78:18:@5303.6]
  wire [3:0] _GEN_202; // @[LoadQueue.scala 76:25:@5289.4]
  wire  _GEN_203; // @[LoadQueue.scala 76:25:@5289.4]
  wire [3:0] _T_2040; // @[:@5311.6]
  wire [3:0] _GEN_205; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_206; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_207; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_208; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_209; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_210; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_211; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_212; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_213; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_214; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_215; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_216; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_217; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_218; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_219; // @[LoadQueue.scala 77:20:@5312.6]
  wire  _GEN_221; // @[LoadQueue.scala 78:18:@5319.6]
  wire  _GEN_222; // @[LoadQueue.scala 78:18:@5319.6]
  wire  _GEN_223; // @[LoadQueue.scala 78:18:@5319.6]
  wire  _GEN_224; // @[LoadQueue.scala 78:18:@5319.6]
  wire  _GEN_225; // @[LoadQueue.scala 78:18:@5319.6]
  wire  _GEN_226; // @[LoadQueue.scala 78:18:@5319.6]
  wire  _GEN_227; // @[LoadQueue.scala 78:18:@5319.6]
  wire  _GEN_228; // @[LoadQueue.scala 78:18:@5319.6]
  wire  _GEN_229; // @[LoadQueue.scala 78:18:@5319.6]
  wire  _GEN_230; // @[LoadQueue.scala 78:18:@5319.6]
  wire  _GEN_231; // @[LoadQueue.scala 78:18:@5319.6]
  wire  _GEN_232; // @[LoadQueue.scala 78:18:@5319.6]
  wire  _GEN_233; // @[LoadQueue.scala 78:18:@5319.6]
  wire  _GEN_234; // @[LoadQueue.scala 78:18:@5319.6]
  wire  _GEN_235; // @[LoadQueue.scala 78:18:@5319.6]
  wire [3:0] _GEN_236; // @[LoadQueue.scala 76:25:@5305.4]
  wire  _GEN_237; // @[LoadQueue.scala 76:25:@5305.4]
  wire [3:0] _T_2058; // @[:@5327.6]
  wire [3:0] _GEN_239; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_240; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_241; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_242; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_243; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_244; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_245; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_246; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_247; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_248; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_249; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_250; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_251; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_252; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_253; // @[LoadQueue.scala 77:20:@5328.6]
  wire  _GEN_255; // @[LoadQueue.scala 78:18:@5335.6]
  wire  _GEN_256; // @[LoadQueue.scala 78:18:@5335.6]
  wire  _GEN_257; // @[LoadQueue.scala 78:18:@5335.6]
  wire  _GEN_258; // @[LoadQueue.scala 78:18:@5335.6]
  wire  _GEN_259; // @[LoadQueue.scala 78:18:@5335.6]
  wire  _GEN_260; // @[LoadQueue.scala 78:18:@5335.6]
  wire  _GEN_261; // @[LoadQueue.scala 78:18:@5335.6]
  wire  _GEN_262; // @[LoadQueue.scala 78:18:@5335.6]
  wire  _GEN_263; // @[LoadQueue.scala 78:18:@5335.6]
  wire  _GEN_264; // @[LoadQueue.scala 78:18:@5335.6]
  wire  _GEN_265; // @[LoadQueue.scala 78:18:@5335.6]
  wire  _GEN_266; // @[LoadQueue.scala 78:18:@5335.6]
  wire  _GEN_267; // @[LoadQueue.scala 78:18:@5335.6]
  wire  _GEN_268; // @[LoadQueue.scala 78:18:@5335.6]
  wire  _GEN_269; // @[LoadQueue.scala 78:18:@5335.6]
  wire [3:0] _GEN_270; // @[LoadQueue.scala 76:25:@5321.4]
  wire  _GEN_271; // @[LoadQueue.scala 76:25:@5321.4]
  wire [3:0] _T_2076; // @[:@5343.6]
  wire [3:0] _GEN_273; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_274; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_275; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_276; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_277; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_278; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_279; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_280; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_281; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_282; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_283; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_284; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_285; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_286; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_287; // @[LoadQueue.scala 77:20:@5344.6]
  wire  _GEN_289; // @[LoadQueue.scala 78:18:@5351.6]
  wire  _GEN_290; // @[LoadQueue.scala 78:18:@5351.6]
  wire  _GEN_291; // @[LoadQueue.scala 78:18:@5351.6]
  wire  _GEN_292; // @[LoadQueue.scala 78:18:@5351.6]
  wire  _GEN_293; // @[LoadQueue.scala 78:18:@5351.6]
  wire  _GEN_294; // @[LoadQueue.scala 78:18:@5351.6]
  wire  _GEN_295; // @[LoadQueue.scala 78:18:@5351.6]
  wire  _GEN_296; // @[LoadQueue.scala 78:18:@5351.6]
  wire  _GEN_297; // @[LoadQueue.scala 78:18:@5351.6]
  wire  _GEN_298; // @[LoadQueue.scala 78:18:@5351.6]
  wire  _GEN_299; // @[LoadQueue.scala 78:18:@5351.6]
  wire  _GEN_300; // @[LoadQueue.scala 78:18:@5351.6]
  wire  _GEN_301; // @[LoadQueue.scala 78:18:@5351.6]
  wire  _GEN_302; // @[LoadQueue.scala 78:18:@5351.6]
  wire  _GEN_303; // @[LoadQueue.scala 78:18:@5351.6]
  wire [3:0] _GEN_304; // @[LoadQueue.scala 76:25:@5337.4]
  wire  _GEN_305; // @[LoadQueue.scala 76:25:@5337.4]
  wire [3:0] _T_2094; // @[:@5359.6]
  wire [3:0] _GEN_307; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_308; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_309; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_310; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_311; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_312; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_313; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_314; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_315; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_316; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_317; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_318; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_319; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_320; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_321; // @[LoadQueue.scala 77:20:@5360.6]
  wire  _GEN_323; // @[LoadQueue.scala 78:18:@5367.6]
  wire  _GEN_324; // @[LoadQueue.scala 78:18:@5367.6]
  wire  _GEN_325; // @[LoadQueue.scala 78:18:@5367.6]
  wire  _GEN_326; // @[LoadQueue.scala 78:18:@5367.6]
  wire  _GEN_327; // @[LoadQueue.scala 78:18:@5367.6]
  wire  _GEN_328; // @[LoadQueue.scala 78:18:@5367.6]
  wire  _GEN_329; // @[LoadQueue.scala 78:18:@5367.6]
  wire  _GEN_330; // @[LoadQueue.scala 78:18:@5367.6]
  wire  _GEN_331; // @[LoadQueue.scala 78:18:@5367.6]
  wire  _GEN_332; // @[LoadQueue.scala 78:18:@5367.6]
  wire  _GEN_333; // @[LoadQueue.scala 78:18:@5367.6]
  wire  _GEN_334; // @[LoadQueue.scala 78:18:@5367.6]
  wire  _GEN_335; // @[LoadQueue.scala 78:18:@5367.6]
  wire  _GEN_336; // @[LoadQueue.scala 78:18:@5367.6]
  wire  _GEN_337; // @[LoadQueue.scala 78:18:@5367.6]
  wire [3:0] _GEN_338; // @[LoadQueue.scala 76:25:@5353.4]
  wire  _GEN_339; // @[LoadQueue.scala 76:25:@5353.4]
  wire [3:0] _T_2112; // @[:@5375.6]
  wire [3:0] _GEN_341; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_342; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_343; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_344; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_345; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_346; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_347; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_348; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_349; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_350; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_351; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_352; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_353; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_354; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_355; // @[LoadQueue.scala 77:20:@5376.6]
  wire  _GEN_357; // @[LoadQueue.scala 78:18:@5383.6]
  wire  _GEN_358; // @[LoadQueue.scala 78:18:@5383.6]
  wire  _GEN_359; // @[LoadQueue.scala 78:18:@5383.6]
  wire  _GEN_360; // @[LoadQueue.scala 78:18:@5383.6]
  wire  _GEN_361; // @[LoadQueue.scala 78:18:@5383.6]
  wire  _GEN_362; // @[LoadQueue.scala 78:18:@5383.6]
  wire  _GEN_363; // @[LoadQueue.scala 78:18:@5383.6]
  wire  _GEN_364; // @[LoadQueue.scala 78:18:@5383.6]
  wire  _GEN_365; // @[LoadQueue.scala 78:18:@5383.6]
  wire  _GEN_366; // @[LoadQueue.scala 78:18:@5383.6]
  wire  _GEN_367; // @[LoadQueue.scala 78:18:@5383.6]
  wire  _GEN_368; // @[LoadQueue.scala 78:18:@5383.6]
  wire  _GEN_369; // @[LoadQueue.scala 78:18:@5383.6]
  wire  _GEN_370; // @[LoadQueue.scala 78:18:@5383.6]
  wire  _GEN_371; // @[LoadQueue.scala 78:18:@5383.6]
  wire [3:0] _GEN_372; // @[LoadQueue.scala 76:25:@5369.4]
  wire  _GEN_373; // @[LoadQueue.scala 76:25:@5369.4]
  wire [3:0] _T_2130; // @[:@5391.6]
  wire [3:0] _GEN_375; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_376; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_377; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_378; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_379; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_380; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_381; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_382; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_383; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_384; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_385; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_386; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_387; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_388; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_389; // @[LoadQueue.scala 77:20:@5392.6]
  wire  _GEN_391; // @[LoadQueue.scala 78:18:@5399.6]
  wire  _GEN_392; // @[LoadQueue.scala 78:18:@5399.6]
  wire  _GEN_393; // @[LoadQueue.scala 78:18:@5399.6]
  wire  _GEN_394; // @[LoadQueue.scala 78:18:@5399.6]
  wire  _GEN_395; // @[LoadQueue.scala 78:18:@5399.6]
  wire  _GEN_396; // @[LoadQueue.scala 78:18:@5399.6]
  wire  _GEN_397; // @[LoadQueue.scala 78:18:@5399.6]
  wire  _GEN_398; // @[LoadQueue.scala 78:18:@5399.6]
  wire  _GEN_399; // @[LoadQueue.scala 78:18:@5399.6]
  wire  _GEN_400; // @[LoadQueue.scala 78:18:@5399.6]
  wire  _GEN_401; // @[LoadQueue.scala 78:18:@5399.6]
  wire  _GEN_402; // @[LoadQueue.scala 78:18:@5399.6]
  wire  _GEN_403; // @[LoadQueue.scala 78:18:@5399.6]
  wire  _GEN_404; // @[LoadQueue.scala 78:18:@5399.6]
  wire  _GEN_405; // @[LoadQueue.scala 78:18:@5399.6]
  wire [3:0] _GEN_406; // @[LoadQueue.scala 76:25:@5385.4]
  wire  _GEN_407; // @[LoadQueue.scala 76:25:@5385.4]
  wire [3:0] _T_2148; // @[:@5407.6]
  wire [3:0] _GEN_409; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_410; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_411; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_412; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_413; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_414; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_415; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_416; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_417; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_418; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_419; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_420; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_421; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_422; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_423; // @[LoadQueue.scala 77:20:@5408.6]
  wire  _GEN_425; // @[LoadQueue.scala 78:18:@5415.6]
  wire  _GEN_426; // @[LoadQueue.scala 78:18:@5415.6]
  wire  _GEN_427; // @[LoadQueue.scala 78:18:@5415.6]
  wire  _GEN_428; // @[LoadQueue.scala 78:18:@5415.6]
  wire  _GEN_429; // @[LoadQueue.scala 78:18:@5415.6]
  wire  _GEN_430; // @[LoadQueue.scala 78:18:@5415.6]
  wire  _GEN_431; // @[LoadQueue.scala 78:18:@5415.6]
  wire  _GEN_432; // @[LoadQueue.scala 78:18:@5415.6]
  wire  _GEN_433; // @[LoadQueue.scala 78:18:@5415.6]
  wire  _GEN_434; // @[LoadQueue.scala 78:18:@5415.6]
  wire  _GEN_435; // @[LoadQueue.scala 78:18:@5415.6]
  wire  _GEN_436; // @[LoadQueue.scala 78:18:@5415.6]
  wire  _GEN_437; // @[LoadQueue.scala 78:18:@5415.6]
  wire  _GEN_438; // @[LoadQueue.scala 78:18:@5415.6]
  wire  _GEN_439; // @[LoadQueue.scala 78:18:@5415.6]
  wire [3:0] _GEN_440; // @[LoadQueue.scala 76:25:@5401.4]
  wire  _GEN_441; // @[LoadQueue.scala 76:25:@5401.4]
  wire [3:0] _T_2166; // @[:@5423.6]
  wire [3:0] _GEN_443; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_444; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_445; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_446; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_447; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_448; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_449; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_450; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_451; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_452; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_453; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_454; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_455; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_456; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_457; // @[LoadQueue.scala 77:20:@5424.6]
  wire  _GEN_459; // @[LoadQueue.scala 78:18:@5431.6]
  wire  _GEN_460; // @[LoadQueue.scala 78:18:@5431.6]
  wire  _GEN_461; // @[LoadQueue.scala 78:18:@5431.6]
  wire  _GEN_462; // @[LoadQueue.scala 78:18:@5431.6]
  wire  _GEN_463; // @[LoadQueue.scala 78:18:@5431.6]
  wire  _GEN_464; // @[LoadQueue.scala 78:18:@5431.6]
  wire  _GEN_465; // @[LoadQueue.scala 78:18:@5431.6]
  wire  _GEN_466; // @[LoadQueue.scala 78:18:@5431.6]
  wire  _GEN_467; // @[LoadQueue.scala 78:18:@5431.6]
  wire  _GEN_468; // @[LoadQueue.scala 78:18:@5431.6]
  wire  _GEN_469; // @[LoadQueue.scala 78:18:@5431.6]
  wire  _GEN_470; // @[LoadQueue.scala 78:18:@5431.6]
  wire  _GEN_471; // @[LoadQueue.scala 78:18:@5431.6]
  wire  _GEN_472; // @[LoadQueue.scala 78:18:@5431.6]
  wire  _GEN_473; // @[LoadQueue.scala 78:18:@5431.6]
  wire [3:0] _GEN_474; // @[LoadQueue.scala 76:25:@5417.4]
  wire  _GEN_475; // @[LoadQueue.scala 76:25:@5417.4]
  wire [3:0] _T_2184; // @[:@5439.6]
  wire [3:0] _GEN_477; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_478; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_479; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_480; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_481; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_482; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_483; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_484; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_485; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_486; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_487; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_488; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_489; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_490; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_491; // @[LoadQueue.scala 77:20:@5440.6]
  wire  _GEN_493; // @[LoadQueue.scala 78:18:@5447.6]
  wire  _GEN_494; // @[LoadQueue.scala 78:18:@5447.6]
  wire  _GEN_495; // @[LoadQueue.scala 78:18:@5447.6]
  wire  _GEN_496; // @[LoadQueue.scala 78:18:@5447.6]
  wire  _GEN_497; // @[LoadQueue.scala 78:18:@5447.6]
  wire  _GEN_498; // @[LoadQueue.scala 78:18:@5447.6]
  wire  _GEN_499; // @[LoadQueue.scala 78:18:@5447.6]
  wire  _GEN_500; // @[LoadQueue.scala 78:18:@5447.6]
  wire  _GEN_501; // @[LoadQueue.scala 78:18:@5447.6]
  wire  _GEN_502; // @[LoadQueue.scala 78:18:@5447.6]
  wire  _GEN_503; // @[LoadQueue.scala 78:18:@5447.6]
  wire  _GEN_504; // @[LoadQueue.scala 78:18:@5447.6]
  wire  _GEN_505; // @[LoadQueue.scala 78:18:@5447.6]
  wire  _GEN_506; // @[LoadQueue.scala 78:18:@5447.6]
  wire  _GEN_507; // @[LoadQueue.scala 78:18:@5447.6]
  wire [3:0] _GEN_508; // @[LoadQueue.scala 76:25:@5433.4]
  wire  _GEN_509; // @[LoadQueue.scala 76:25:@5433.4]
  wire [3:0] _T_2202; // @[:@5455.6]
  wire [3:0] _GEN_511; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_512; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_513; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_514; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_515; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_516; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_517; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_518; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_519; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_520; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_521; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_522; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_523; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_524; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_525; // @[LoadQueue.scala 77:20:@5456.6]
  wire  _GEN_527; // @[LoadQueue.scala 78:18:@5463.6]
  wire  _GEN_528; // @[LoadQueue.scala 78:18:@5463.6]
  wire  _GEN_529; // @[LoadQueue.scala 78:18:@5463.6]
  wire  _GEN_530; // @[LoadQueue.scala 78:18:@5463.6]
  wire  _GEN_531; // @[LoadQueue.scala 78:18:@5463.6]
  wire  _GEN_532; // @[LoadQueue.scala 78:18:@5463.6]
  wire  _GEN_533; // @[LoadQueue.scala 78:18:@5463.6]
  wire  _GEN_534; // @[LoadQueue.scala 78:18:@5463.6]
  wire  _GEN_535; // @[LoadQueue.scala 78:18:@5463.6]
  wire  _GEN_536; // @[LoadQueue.scala 78:18:@5463.6]
  wire  _GEN_537; // @[LoadQueue.scala 78:18:@5463.6]
  wire  _GEN_538; // @[LoadQueue.scala 78:18:@5463.6]
  wire  _GEN_539; // @[LoadQueue.scala 78:18:@5463.6]
  wire  _GEN_540; // @[LoadQueue.scala 78:18:@5463.6]
  wire  _GEN_541; // @[LoadQueue.scala 78:18:@5463.6]
  wire [3:0] _GEN_542; // @[LoadQueue.scala 76:25:@5449.4]
  wire  _GEN_543; // @[LoadQueue.scala 76:25:@5449.4]
  reg [3:0] previousStoreHead; // @[LoadQueue.scala 93:34:@5465.4]
  reg [31:0] _RAND_162;
  wire [4:0] _T_2224; // @[util.scala 10:8:@5474.6]
  wire [4:0] _GEN_272; // @[util.scala 10:14:@5475.6]
  wire [4:0] _T_2225; // @[util.scala 10:14:@5475.6]
  wire [4:0] _GEN_2377; // @[LoadQueue.scala 97:56:@5476.6]
  wire  _T_2226; // @[LoadQueue.scala 97:56:@5476.6]
  wire  _T_2227; // @[LoadQueue.scala 96:50:@5477.6]
  wire  _T_2229; // @[LoadQueue.scala 96:34:@5478.6]
  wire  _T_2231; // @[LoadQueue.scala 101:36:@5486.8]
  wire  _T_2232; // @[LoadQueue.scala 101:86:@5487.8]
  wire  _T_2233; // @[LoadQueue.scala 101:61:@5488.8]
  wire  _T_2235; // @[LoadQueue.scala 103:36:@5493.10]
  wire  _T_2236; // @[LoadQueue.scala 103:69:@5494.10]
  wire  _T_2237; // @[LoadQueue.scala 104:31:@5495.10]
  wire  _T_2238; // @[LoadQueue.scala 103:94:@5496.10]
  wire  _T_2240; // @[LoadQueue.scala 103:54:@5497.10]
  wire  _T_2241; // @[LoadQueue.scala 103:51:@5498.10]
  wire  _GEN_560; // @[LoadQueue.scala 104:53:@5499.10]
  wire  _GEN_561; // @[LoadQueue.scala 101:102:@5489.8]
  wire  _GEN_562; // @[LoadQueue.scala 99:27:@5482.6]
  wire  _GEN_563; // @[LoadQueue.scala 95:34:@5467.4]
  wire [4:0] _T_2254; // @[util.scala 10:8:@5510.6]
  wire [4:0] _GEN_288; // @[util.scala 10:14:@5511.6]
  wire [4:0] _T_2255; // @[util.scala 10:14:@5511.6]
  wire  _T_2256; // @[LoadQueue.scala 97:56:@5512.6]
  wire  _T_2257; // @[LoadQueue.scala 96:50:@5513.6]
  wire  _T_2259; // @[LoadQueue.scala 96:34:@5514.6]
  wire  _T_2261; // @[LoadQueue.scala 101:36:@5522.8]
  wire  _T_2262; // @[LoadQueue.scala 101:86:@5523.8]
  wire  _T_2263; // @[LoadQueue.scala 101:61:@5524.8]
  wire  _T_2266; // @[LoadQueue.scala 103:69:@5530.10]
  wire  _T_2267; // @[LoadQueue.scala 104:31:@5531.10]
  wire  _T_2268; // @[LoadQueue.scala 103:94:@5532.10]
  wire  _T_2270; // @[LoadQueue.scala 103:54:@5533.10]
  wire  _T_2271; // @[LoadQueue.scala 103:51:@5534.10]
  wire  _GEN_580; // @[LoadQueue.scala 104:53:@5535.10]
  wire  _GEN_581; // @[LoadQueue.scala 101:102:@5525.8]
  wire  _GEN_582; // @[LoadQueue.scala 99:27:@5518.6]
  wire  _GEN_583; // @[LoadQueue.scala 95:34:@5503.4]
  wire [4:0] _T_2284; // @[util.scala 10:8:@5546.6]
  wire [4:0] _GEN_306; // @[util.scala 10:14:@5547.6]
  wire [4:0] _T_2285; // @[util.scala 10:14:@5547.6]
  wire  _T_2286; // @[LoadQueue.scala 97:56:@5548.6]
  wire  _T_2287; // @[LoadQueue.scala 96:50:@5549.6]
  wire  _T_2289; // @[LoadQueue.scala 96:34:@5550.6]
  wire  _T_2291; // @[LoadQueue.scala 101:36:@5558.8]
  wire  _T_2292; // @[LoadQueue.scala 101:86:@5559.8]
  wire  _T_2293; // @[LoadQueue.scala 101:61:@5560.8]
  wire  _T_2296; // @[LoadQueue.scala 103:69:@5566.10]
  wire  _T_2297; // @[LoadQueue.scala 104:31:@5567.10]
  wire  _T_2298; // @[LoadQueue.scala 103:94:@5568.10]
  wire  _T_2300; // @[LoadQueue.scala 103:54:@5569.10]
  wire  _T_2301; // @[LoadQueue.scala 103:51:@5570.10]
  wire  _GEN_600; // @[LoadQueue.scala 104:53:@5571.10]
  wire  _GEN_601; // @[LoadQueue.scala 101:102:@5561.8]
  wire  _GEN_602; // @[LoadQueue.scala 99:27:@5554.6]
  wire  _GEN_603; // @[LoadQueue.scala 95:34:@5539.4]
  wire [4:0] _T_2314; // @[util.scala 10:8:@5582.6]
  wire [4:0] _GEN_322; // @[util.scala 10:14:@5583.6]
  wire [4:0] _T_2315; // @[util.scala 10:14:@5583.6]
  wire  _T_2316; // @[LoadQueue.scala 97:56:@5584.6]
  wire  _T_2317; // @[LoadQueue.scala 96:50:@5585.6]
  wire  _T_2319; // @[LoadQueue.scala 96:34:@5586.6]
  wire  _T_2321; // @[LoadQueue.scala 101:36:@5594.8]
  wire  _T_2322; // @[LoadQueue.scala 101:86:@5595.8]
  wire  _T_2323; // @[LoadQueue.scala 101:61:@5596.8]
  wire  _T_2326; // @[LoadQueue.scala 103:69:@5602.10]
  wire  _T_2327; // @[LoadQueue.scala 104:31:@5603.10]
  wire  _T_2328; // @[LoadQueue.scala 103:94:@5604.10]
  wire  _T_2330; // @[LoadQueue.scala 103:54:@5605.10]
  wire  _T_2331; // @[LoadQueue.scala 103:51:@5606.10]
  wire  _GEN_620; // @[LoadQueue.scala 104:53:@5607.10]
  wire  _GEN_621; // @[LoadQueue.scala 101:102:@5597.8]
  wire  _GEN_622; // @[LoadQueue.scala 99:27:@5590.6]
  wire  _GEN_623; // @[LoadQueue.scala 95:34:@5575.4]
  wire [4:0] _T_2344; // @[util.scala 10:8:@5618.6]
  wire [4:0] _GEN_340; // @[util.scala 10:14:@5619.6]
  wire [4:0] _T_2345; // @[util.scala 10:14:@5619.6]
  wire  _T_2346; // @[LoadQueue.scala 97:56:@5620.6]
  wire  _T_2347; // @[LoadQueue.scala 96:50:@5621.6]
  wire  _T_2349; // @[LoadQueue.scala 96:34:@5622.6]
  wire  _T_2351; // @[LoadQueue.scala 101:36:@5630.8]
  wire  _T_2352; // @[LoadQueue.scala 101:86:@5631.8]
  wire  _T_2353; // @[LoadQueue.scala 101:61:@5632.8]
  wire  _T_2356; // @[LoadQueue.scala 103:69:@5638.10]
  wire  _T_2357; // @[LoadQueue.scala 104:31:@5639.10]
  wire  _T_2358; // @[LoadQueue.scala 103:94:@5640.10]
  wire  _T_2360; // @[LoadQueue.scala 103:54:@5641.10]
  wire  _T_2361; // @[LoadQueue.scala 103:51:@5642.10]
  wire  _GEN_640; // @[LoadQueue.scala 104:53:@5643.10]
  wire  _GEN_641; // @[LoadQueue.scala 101:102:@5633.8]
  wire  _GEN_642; // @[LoadQueue.scala 99:27:@5626.6]
  wire  _GEN_643; // @[LoadQueue.scala 95:34:@5611.4]
  wire [4:0] _T_2374; // @[util.scala 10:8:@5654.6]
  wire [4:0] _GEN_356; // @[util.scala 10:14:@5655.6]
  wire [4:0] _T_2375; // @[util.scala 10:14:@5655.6]
  wire  _T_2376; // @[LoadQueue.scala 97:56:@5656.6]
  wire  _T_2377; // @[LoadQueue.scala 96:50:@5657.6]
  wire  _T_2379; // @[LoadQueue.scala 96:34:@5658.6]
  wire  _T_2381; // @[LoadQueue.scala 101:36:@5666.8]
  wire  _T_2382; // @[LoadQueue.scala 101:86:@5667.8]
  wire  _T_2383; // @[LoadQueue.scala 101:61:@5668.8]
  wire  _T_2386; // @[LoadQueue.scala 103:69:@5674.10]
  wire  _T_2387; // @[LoadQueue.scala 104:31:@5675.10]
  wire  _T_2388; // @[LoadQueue.scala 103:94:@5676.10]
  wire  _T_2390; // @[LoadQueue.scala 103:54:@5677.10]
  wire  _T_2391; // @[LoadQueue.scala 103:51:@5678.10]
  wire  _GEN_660; // @[LoadQueue.scala 104:53:@5679.10]
  wire  _GEN_661; // @[LoadQueue.scala 101:102:@5669.8]
  wire  _GEN_662; // @[LoadQueue.scala 99:27:@5662.6]
  wire  _GEN_663; // @[LoadQueue.scala 95:34:@5647.4]
  wire [4:0] _T_2404; // @[util.scala 10:8:@5690.6]
  wire [4:0] _GEN_374; // @[util.scala 10:14:@5691.6]
  wire [4:0] _T_2405; // @[util.scala 10:14:@5691.6]
  wire  _T_2406; // @[LoadQueue.scala 97:56:@5692.6]
  wire  _T_2407; // @[LoadQueue.scala 96:50:@5693.6]
  wire  _T_2409; // @[LoadQueue.scala 96:34:@5694.6]
  wire  _T_2411; // @[LoadQueue.scala 101:36:@5702.8]
  wire  _T_2412; // @[LoadQueue.scala 101:86:@5703.8]
  wire  _T_2413; // @[LoadQueue.scala 101:61:@5704.8]
  wire  _T_2416; // @[LoadQueue.scala 103:69:@5710.10]
  wire  _T_2417; // @[LoadQueue.scala 104:31:@5711.10]
  wire  _T_2418; // @[LoadQueue.scala 103:94:@5712.10]
  wire  _T_2420; // @[LoadQueue.scala 103:54:@5713.10]
  wire  _T_2421; // @[LoadQueue.scala 103:51:@5714.10]
  wire  _GEN_680; // @[LoadQueue.scala 104:53:@5715.10]
  wire  _GEN_681; // @[LoadQueue.scala 101:102:@5705.8]
  wire  _GEN_682; // @[LoadQueue.scala 99:27:@5698.6]
  wire  _GEN_683; // @[LoadQueue.scala 95:34:@5683.4]
  wire [4:0] _T_2434; // @[util.scala 10:8:@5726.6]
  wire [4:0] _GEN_390; // @[util.scala 10:14:@5727.6]
  wire [4:0] _T_2435; // @[util.scala 10:14:@5727.6]
  wire  _T_2436; // @[LoadQueue.scala 97:56:@5728.6]
  wire  _T_2437; // @[LoadQueue.scala 96:50:@5729.6]
  wire  _T_2439; // @[LoadQueue.scala 96:34:@5730.6]
  wire  _T_2441; // @[LoadQueue.scala 101:36:@5738.8]
  wire  _T_2442; // @[LoadQueue.scala 101:86:@5739.8]
  wire  _T_2443; // @[LoadQueue.scala 101:61:@5740.8]
  wire  _T_2446; // @[LoadQueue.scala 103:69:@5746.10]
  wire  _T_2447; // @[LoadQueue.scala 104:31:@5747.10]
  wire  _T_2448; // @[LoadQueue.scala 103:94:@5748.10]
  wire  _T_2450; // @[LoadQueue.scala 103:54:@5749.10]
  wire  _T_2451; // @[LoadQueue.scala 103:51:@5750.10]
  wire  _GEN_700; // @[LoadQueue.scala 104:53:@5751.10]
  wire  _GEN_701; // @[LoadQueue.scala 101:102:@5741.8]
  wire  _GEN_702; // @[LoadQueue.scala 99:27:@5734.6]
  wire  _GEN_703; // @[LoadQueue.scala 95:34:@5719.4]
  wire [4:0] _T_2464; // @[util.scala 10:8:@5762.6]
  wire [4:0] _GEN_408; // @[util.scala 10:14:@5763.6]
  wire [4:0] _T_2465; // @[util.scala 10:14:@5763.6]
  wire  _T_2466; // @[LoadQueue.scala 97:56:@5764.6]
  wire  _T_2467; // @[LoadQueue.scala 96:50:@5765.6]
  wire  _T_2469; // @[LoadQueue.scala 96:34:@5766.6]
  wire  _T_2471; // @[LoadQueue.scala 101:36:@5774.8]
  wire  _T_2472; // @[LoadQueue.scala 101:86:@5775.8]
  wire  _T_2473; // @[LoadQueue.scala 101:61:@5776.8]
  wire  _T_2476; // @[LoadQueue.scala 103:69:@5782.10]
  wire  _T_2477; // @[LoadQueue.scala 104:31:@5783.10]
  wire  _T_2478; // @[LoadQueue.scala 103:94:@5784.10]
  wire  _T_2480; // @[LoadQueue.scala 103:54:@5785.10]
  wire  _T_2481; // @[LoadQueue.scala 103:51:@5786.10]
  wire  _GEN_720; // @[LoadQueue.scala 104:53:@5787.10]
  wire  _GEN_721; // @[LoadQueue.scala 101:102:@5777.8]
  wire  _GEN_722; // @[LoadQueue.scala 99:27:@5770.6]
  wire  _GEN_723; // @[LoadQueue.scala 95:34:@5755.4]
  wire [4:0] _T_2494; // @[util.scala 10:8:@5798.6]
  wire [4:0] _GEN_424; // @[util.scala 10:14:@5799.6]
  wire [4:0] _T_2495; // @[util.scala 10:14:@5799.6]
  wire  _T_2496; // @[LoadQueue.scala 97:56:@5800.6]
  wire  _T_2497; // @[LoadQueue.scala 96:50:@5801.6]
  wire  _T_2499; // @[LoadQueue.scala 96:34:@5802.6]
  wire  _T_2501; // @[LoadQueue.scala 101:36:@5810.8]
  wire  _T_2502; // @[LoadQueue.scala 101:86:@5811.8]
  wire  _T_2503; // @[LoadQueue.scala 101:61:@5812.8]
  wire  _T_2506; // @[LoadQueue.scala 103:69:@5818.10]
  wire  _T_2507; // @[LoadQueue.scala 104:31:@5819.10]
  wire  _T_2508; // @[LoadQueue.scala 103:94:@5820.10]
  wire  _T_2510; // @[LoadQueue.scala 103:54:@5821.10]
  wire  _T_2511; // @[LoadQueue.scala 103:51:@5822.10]
  wire  _GEN_740; // @[LoadQueue.scala 104:53:@5823.10]
  wire  _GEN_741; // @[LoadQueue.scala 101:102:@5813.8]
  wire  _GEN_742; // @[LoadQueue.scala 99:27:@5806.6]
  wire  _GEN_743; // @[LoadQueue.scala 95:34:@5791.4]
  wire [4:0] _T_2524; // @[util.scala 10:8:@5834.6]
  wire [4:0] _GEN_442; // @[util.scala 10:14:@5835.6]
  wire [4:0] _T_2525; // @[util.scala 10:14:@5835.6]
  wire  _T_2526; // @[LoadQueue.scala 97:56:@5836.6]
  wire  _T_2527; // @[LoadQueue.scala 96:50:@5837.6]
  wire  _T_2529; // @[LoadQueue.scala 96:34:@5838.6]
  wire  _T_2531; // @[LoadQueue.scala 101:36:@5846.8]
  wire  _T_2532; // @[LoadQueue.scala 101:86:@5847.8]
  wire  _T_2533; // @[LoadQueue.scala 101:61:@5848.8]
  wire  _T_2536; // @[LoadQueue.scala 103:69:@5854.10]
  wire  _T_2537; // @[LoadQueue.scala 104:31:@5855.10]
  wire  _T_2538; // @[LoadQueue.scala 103:94:@5856.10]
  wire  _T_2540; // @[LoadQueue.scala 103:54:@5857.10]
  wire  _T_2541; // @[LoadQueue.scala 103:51:@5858.10]
  wire  _GEN_760; // @[LoadQueue.scala 104:53:@5859.10]
  wire  _GEN_761; // @[LoadQueue.scala 101:102:@5849.8]
  wire  _GEN_762; // @[LoadQueue.scala 99:27:@5842.6]
  wire  _GEN_763; // @[LoadQueue.scala 95:34:@5827.4]
  wire [4:0] _T_2554; // @[util.scala 10:8:@5870.6]
  wire [4:0] _GEN_458; // @[util.scala 10:14:@5871.6]
  wire [4:0] _T_2555; // @[util.scala 10:14:@5871.6]
  wire  _T_2556; // @[LoadQueue.scala 97:56:@5872.6]
  wire  _T_2557; // @[LoadQueue.scala 96:50:@5873.6]
  wire  _T_2559; // @[LoadQueue.scala 96:34:@5874.6]
  wire  _T_2561; // @[LoadQueue.scala 101:36:@5882.8]
  wire  _T_2562; // @[LoadQueue.scala 101:86:@5883.8]
  wire  _T_2563; // @[LoadQueue.scala 101:61:@5884.8]
  wire  _T_2566; // @[LoadQueue.scala 103:69:@5890.10]
  wire  _T_2567; // @[LoadQueue.scala 104:31:@5891.10]
  wire  _T_2568; // @[LoadQueue.scala 103:94:@5892.10]
  wire  _T_2570; // @[LoadQueue.scala 103:54:@5893.10]
  wire  _T_2571; // @[LoadQueue.scala 103:51:@5894.10]
  wire  _GEN_780; // @[LoadQueue.scala 104:53:@5895.10]
  wire  _GEN_781; // @[LoadQueue.scala 101:102:@5885.8]
  wire  _GEN_782; // @[LoadQueue.scala 99:27:@5878.6]
  wire  _GEN_783; // @[LoadQueue.scala 95:34:@5863.4]
  wire [4:0] _T_2584; // @[util.scala 10:8:@5906.6]
  wire [4:0] _GEN_476; // @[util.scala 10:14:@5907.6]
  wire [4:0] _T_2585; // @[util.scala 10:14:@5907.6]
  wire  _T_2586; // @[LoadQueue.scala 97:56:@5908.6]
  wire  _T_2587; // @[LoadQueue.scala 96:50:@5909.6]
  wire  _T_2589; // @[LoadQueue.scala 96:34:@5910.6]
  wire  _T_2591; // @[LoadQueue.scala 101:36:@5918.8]
  wire  _T_2592; // @[LoadQueue.scala 101:86:@5919.8]
  wire  _T_2593; // @[LoadQueue.scala 101:61:@5920.8]
  wire  _T_2596; // @[LoadQueue.scala 103:69:@5926.10]
  wire  _T_2597; // @[LoadQueue.scala 104:31:@5927.10]
  wire  _T_2598; // @[LoadQueue.scala 103:94:@5928.10]
  wire  _T_2600; // @[LoadQueue.scala 103:54:@5929.10]
  wire  _T_2601; // @[LoadQueue.scala 103:51:@5930.10]
  wire  _GEN_800; // @[LoadQueue.scala 104:53:@5931.10]
  wire  _GEN_801; // @[LoadQueue.scala 101:102:@5921.8]
  wire  _GEN_802; // @[LoadQueue.scala 99:27:@5914.6]
  wire  _GEN_803; // @[LoadQueue.scala 95:34:@5899.4]
  wire [4:0] _T_2614; // @[util.scala 10:8:@5942.6]
  wire [4:0] _GEN_492; // @[util.scala 10:14:@5943.6]
  wire [4:0] _T_2615; // @[util.scala 10:14:@5943.6]
  wire  _T_2616; // @[LoadQueue.scala 97:56:@5944.6]
  wire  _T_2617; // @[LoadQueue.scala 96:50:@5945.6]
  wire  _T_2619; // @[LoadQueue.scala 96:34:@5946.6]
  wire  _T_2621; // @[LoadQueue.scala 101:36:@5954.8]
  wire  _T_2622; // @[LoadQueue.scala 101:86:@5955.8]
  wire  _T_2623; // @[LoadQueue.scala 101:61:@5956.8]
  wire  _T_2626; // @[LoadQueue.scala 103:69:@5962.10]
  wire  _T_2627; // @[LoadQueue.scala 104:31:@5963.10]
  wire  _T_2628; // @[LoadQueue.scala 103:94:@5964.10]
  wire  _T_2630; // @[LoadQueue.scala 103:54:@5965.10]
  wire  _T_2631; // @[LoadQueue.scala 103:51:@5966.10]
  wire  _GEN_820; // @[LoadQueue.scala 104:53:@5967.10]
  wire  _GEN_821; // @[LoadQueue.scala 101:102:@5957.8]
  wire  _GEN_822; // @[LoadQueue.scala 99:27:@5950.6]
  wire  _GEN_823; // @[LoadQueue.scala 95:34:@5935.4]
  wire [4:0] _T_2644; // @[util.scala 10:8:@5978.6]
  wire [4:0] _GEN_510; // @[util.scala 10:14:@5979.6]
  wire [4:0] _T_2645; // @[util.scala 10:14:@5979.6]
  wire  _T_2646; // @[LoadQueue.scala 97:56:@5980.6]
  wire  _T_2647; // @[LoadQueue.scala 96:50:@5981.6]
  wire  _T_2649; // @[LoadQueue.scala 96:34:@5982.6]
  wire  _T_2651; // @[LoadQueue.scala 101:36:@5990.8]
  wire  _T_2652; // @[LoadQueue.scala 101:86:@5991.8]
  wire  _T_2653; // @[LoadQueue.scala 101:61:@5992.8]
  wire  _T_2656; // @[LoadQueue.scala 103:69:@5998.10]
  wire  _T_2657; // @[LoadQueue.scala 104:31:@5999.10]
  wire  _T_2658; // @[LoadQueue.scala 103:94:@6000.10]
  wire  _T_2660; // @[LoadQueue.scala 103:54:@6001.10]
  wire  _T_2661; // @[LoadQueue.scala 103:51:@6002.10]
  wire  _GEN_840; // @[LoadQueue.scala 104:53:@6003.10]
  wire  _GEN_841; // @[LoadQueue.scala 101:102:@5993.8]
  wire  _GEN_842; // @[LoadQueue.scala 99:27:@5986.6]
  wire  _GEN_843; // @[LoadQueue.scala 95:34:@5971.4]
  wire [4:0] _T_2674; // @[util.scala 10:8:@6014.6]
  wire [4:0] _GEN_526; // @[util.scala 10:14:@6015.6]
  wire [4:0] _T_2675; // @[util.scala 10:14:@6015.6]
  wire  _T_2676; // @[LoadQueue.scala 97:56:@6016.6]
  wire  _T_2677; // @[LoadQueue.scala 96:50:@6017.6]
  wire  _T_2679; // @[LoadQueue.scala 96:34:@6018.6]
  wire  _T_2681; // @[LoadQueue.scala 101:36:@6026.8]
  wire  _T_2682; // @[LoadQueue.scala 101:86:@6027.8]
  wire  _T_2683; // @[LoadQueue.scala 101:61:@6028.8]
  wire  _T_2686; // @[LoadQueue.scala 103:69:@6034.10]
  wire  _T_2687; // @[LoadQueue.scala 104:31:@6035.10]
  wire  _T_2688; // @[LoadQueue.scala 103:94:@6036.10]
  wire  _T_2690; // @[LoadQueue.scala 103:54:@6037.10]
  wire  _T_2691; // @[LoadQueue.scala 103:51:@6038.10]
  wire  _GEN_860; // @[LoadQueue.scala 104:53:@6039.10]
  wire  _GEN_861; // @[LoadQueue.scala 101:102:@6029.8]
  wire  _GEN_862; // @[LoadQueue.scala 99:27:@6022.6]
  wire  _GEN_863; // @[LoadQueue.scala 95:34:@6007.4]
  wire [15:0] _T_2695; // @[OneHot.scala 52:12:@6044.4]
  wire  _T_2697; // @[util.scala 60:60:@6046.4]
  wire  _T_2698; // @[util.scala 60:60:@6047.4]
  wire  _T_2699; // @[util.scala 60:60:@6048.4]
  wire  _T_2700; // @[util.scala 60:60:@6049.4]
  wire  _T_2701; // @[util.scala 60:60:@6050.4]
  wire  _T_2702; // @[util.scala 60:60:@6051.4]
  wire  _T_2703; // @[util.scala 60:60:@6052.4]
  wire  _T_2704; // @[util.scala 60:60:@6053.4]
  wire  _T_2705; // @[util.scala 60:60:@6054.4]
  wire  _T_2706; // @[util.scala 60:60:@6055.4]
  wire  _T_2707; // @[util.scala 60:60:@6056.4]
  wire  _T_2708; // @[util.scala 60:60:@6057.4]
  wire  _T_2709; // @[util.scala 60:60:@6058.4]
  wire  _T_2710; // @[util.scala 60:60:@6059.4]
  wire  _T_2711; // @[util.scala 60:60:@6060.4]
  wire  _T_2712; // @[util.scala 60:60:@6061.4]
  wire [255:0] _T_4843; // @[Mux.scala 19:72:@7585.4]
  wire [255:0] _T_4850; // @[Mux.scala 19:72:@7592.4]
  wire [511:0] _T_4851; // @[Mux.scala 19:72:@7593.4]
  wire [511:0] _T_4853; // @[Mux.scala 19:72:@7594.4]
  wire [255:0] _T_4860; // @[Mux.scala 19:72:@7601.4]
  wire [255:0] _T_4867; // @[Mux.scala 19:72:@7608.4]
  wire [511:0] _T_4868; // @[Mux.scala 19:72:@7609.4]
  wire [511:0] _T_4870; // @[Mux.scala 19:72:@7610.4]
  wire [255:0] _T_4877; // @[Mux.scala 19:72:@7617.4]
  wire [255:0] _T_4884; // @[Mux.scala 19:72:@7624.4]
  wire [511:0] _T_4885; // @[Mux.scala 19:72:@7625.4]
  wire [511:0] _T_4887; // @[Mux.scala 19:72:@7626.4]
  wire [255:0] _T_4894; // @[Mux.scala 19:72:@7633.4]
  wire [255:0] _T_4901; // @[Mux.scala 19:72:@7640.4]
  wire [511:0] _T_4902; // @[Mux.scala 19:72:@7641.4]
  wire [511:0] _T_4904; // @[Mux.scala 19:72:@7642.4]
  wire [255:0] _T_4911; // @[Mux.scala 19:72:@7649.4]
  wire [255:0] _T_4918; // @[Mux.scala 19:72:@7656.4]
  wire [511:0] _T_4919; // @[Mux.scala 19:72:@7657.4]
  wire [511:0] _T_4921; // @[Mux.scala 19:72:@7658.4]
  wire [255:0] _T_4928; // @[Mux.scala 19:72:@7665.4]
  wire [255:0] _T_4935; // @[Mux.scala 19:72:@7672.4]
  wire [511:0] _T_4936; // @[Mux.scala 19:72:@7673.4]
  wire [511:0] _T_4938; // @[Mux.scala 19:72:@7674.4]
  wire [255:0] _T_4945; // @[Mux.scala 19:72:@7681.4]
  wire [255:0] _T_4952; // @[Mux.scala 19:72:@7688.4]
  wire [511:0] _T_4953; // @[Mux.scala 19:72:@7689.4]
  wire [511:0] _T_4955; // @[Mux.scala 19:72:@7690.4]
  wire [255:0] _T_4962; // @[Mux.scala 19:72:@7697.4]
  wire [255:0] _T_4969; // @[Mux.scala 19:72:@7704.4]
  wire [511:0] _T_4970; // @[Mux.scala 19:72:@7705.4]
  wire [511:0] _T_4972; // @[Mux.scala 19:72:@7706.4]
  wire [511:0] _T_4987; // @[Mux.scala 19:72:@7721.4]
  wire [511:0] _T_4989; // @[Mux.scala 19:72:@7722.4]
  wire [511:0] _T_5004; // @[Mux.scala 19:72:@7737.4]
  wire [511:0] _T_5006; // @[Mux.scala 19:72:@7738.4]
  wire [511:0] _T_5021; // @[Mux.scala 19:72:@7753.4]
  wire [511:0] _T_5023; // @[Mux.scala 19:72:@7754.4]
  wire [511:0] _T_5038; // @[Mux.scala 19:72:@7769.4]
  wire [511:0] _T_5040; // @[Mux.scala 19:72:@7770.4]
  wire [511:0] _T_5055; // @[Mux.scala 19:72:@7785.4]
  wire [511:0] _T_5057; // @[Mux.scala 19:72:@7786.4]
  wire [511:0] _T_5072; // @[Mux.scala 19:72:@7801.4]
  wire [511:0] _T_5074; // @[Mux.scala 19:72:@7802.4]
  wire [511:0] _T_5089; // @[Mux.scala 19:72:@7817.4]
  wire [511:0] _T_5091; // @[Mux.scala 19:72:@7818.4]
  wire [511:0] _T_5106; // @[Mux.scala 19:72:@7833.4]
  wire [511:0] _T_5108; // @[Mux.scala 19:72:@7834.4]
  wire [511:0] _T_5109; // @[Mux.scala 19:72:@7835.4]
  wire [511:0] _T_5110; // @[Mux.scala 19:72:@7836.4]
  wire [511:0] _T_5111; // @[Mux.scala 19:72:@7837.4]
  wire [511:0] _T_5112; // @[Mux.scala 19:72:@7838.4]
  wire [511:0] _T_5113; // @[Mux.scala 19:72:@7839.4]
  wire [511:0] _T_5114; // @[Mux.scala 19:72:@7840.4]
  wire [511:0] _T_5115; // @[Mux.scala 19:72:@7841.4]
  wire [511:0] _T_5116; // @[Mux.scala 19:72:@7842.4]
  wire [511:0] _T_5117; // @[Mux.scala 19:72:@7843.4]
  wire [511:0] _T_5118; // @[Mux.scala 19:72:@7844.4]
  wire [511:0] _T_5119; // @[Mux.scala 19:72:@7845.4]
  wire [511:0] _T_5120; // @[Mux.scala 19:72:@7846.4]
  wire [511:0] _T_5121; // @[Mux.scala 19:72:@7847.4]
  wire [511:0] _T_5122; // @[Mux.scala 19:72:@7848.4]
  wire [511:0] _T_5123; // @[Mux.scala 19:72:@7849.4]
  wire [7:0] _T_5700; // @[Mux.scala 19:72:@8199.4]
  wire [7:0] _T_5707; // @[Mux.scala 19:72:@8206.4]
  wire [15:0] _T_5708; // @[Mux.scala 19:72:@8207.4]
  wire [15:0] _T_5710; // @[Mux.scala 19:72:@8208.4]
  wire [7:0] _T_5717; // @[Mux.scala 19:72:@8215.4]
  wire [7:0] _T_5724; // @[Mux.scala 19:72:@8222.4]
  wire [15:0] _T_5725; // @[Mux.scala 19:72:@8223.4]
  wire [15:0] _T_5727; // @[Mux.scala 19:72:@8224.4]
  wire [7:0] _T_5734; // @[Mux.scala 19:72:@8231.4]
  wire [7:0] _T_5741; // @[Mux.scala 19:72:@8238.4]
  wire [15:0] _T_5742; // @[Mux.scala 19:72:@8239.4]
  wire [15:0] _T_5744; // @[Mux.scala 19:72:@8240.4]
  wire [7:0] _T_5751; // @[Mux.scala 19:72:@8247.4]
  wire [7:0] _T_5758; // @[Mux.scala 19:72:@8254.4]
  wire [15:0] _T_5759; // @[Mux.scala 19:72:@8255.4]
  wire [15:0] _T_5761; // @[Mux.scala 19:72:@8256.4]
  wire [7:0] _T_5768; // @[Mux.scala 19:72:@8263.4]
  wire [7:0] _T_5775; // @[Mux.scala 19:72:@8270.4]
  wire [15:0] _T_5776; // @[Mux.scala 19:72:@8271.4]
  wire [15:0] _T_5778; // @[Mux.scala 19:72:@8272.4]
  wire [7:0] _T_5785; // @[Mux.scala 19:72:@8279.4]
  wire [7:0] _T_5792; // @[Mux.scala 19:72:@8286.4]
  wire [15:0] _T_5793; // @[Mux.scala 19:72:@8287.4]
  wire [15:0] _T_5795; // @[Mux.scala 19:72:@8288.4]
  wire [7:0] _T_5802; // @[Mux.scala 19:72:@8295.4]
  wire [7:0] _T_5809; // @[Mux.scala 19:72:@8302.4]
  wire [15:0] _T_5810; // @[Mux.scala 19:72:@8303.4]
  wire [15:0] _T_5812; // @[Mux.scala 19:72:@8304.4]
  wire [7:0] _T_5819; // @[Mux.scala 19:72:@8311.4]
  wire [7:0] _T_5826; // @[Mux.scala 19:72:@8318.4]
  wire [15:0] _T_5827; // @[Mux.scala 19:72:@8319.4]
  wire [15:0] _T_5829; // @[Mux.scala 19:72:@8320.4]
  wire [15:0] _T_5844; // @[Mux.scala 19:72:@8335.4]
  wire [15:0] _T_5846; // @[Mux.scala 19:72:@8336.4]
  wire [15:0] _T_5861; // @[Mux.scala 19:72:@8351.4]
  wire [15:0] _T_5863; // @[Mux.scala 19:72:@8352.4]
  wire [15:0] _T_5878; // @[Mux.scala 19:72:@8367.4]
  wire [15:0] _T_5880; // @[Mux.scala 19:72:@8368.4]
  wire [15:0] _T_5895; // @[Mux.scala 19:72:@8383.4]
  wire [15:0] _T_5897; // @[Mux.scala 19:72:@8384.4]
  wire [15:0] _T_5912; // @[Mux.scala 19:72:@8399.4]
  wire [15:0] _T_5914; // @[Mux.scala 19:72:@8400.4]
  wire [15:0] _T_5929; // @[Mux.scala 19:72:@8415.4]
  wire [15:0] _T_5931; // @[Mux.scala 19:72:@8416.4]
  wire [15:0] _T_5946; // @[Mux.scala 19:72:@8431.4]
  wire [15:0] _T_5948; // @[Mux.scala 19:72:@8432.4]
  wire [15:0] _T_5963; // @[Mux.scala 19:72:@8447.4]
  wire [15:0] _T_5965; // @[Mux.scala 19:72:@8448.4]
  wire [15:0] _T_5966; // @[Mux.scala 19:72:@8449.4]
  wire [15:0] _T_5967; // @[Mux.scala 19:72:@8450.4]
  wire [15:0] _T_5968; // @[Mux.scala 19:72:@8451.4]
  wire [15:0] _T_5969; // @[Mux.scala 19:72:@8452.4]
  wire [15:0] _T_5970; // @[Mux.scala 19:72:@8453.4]
  wire [15:0] _T_5971; // @[Mux.scala 19:72:@8454.4]
  wire [15:0] _T_5972; // @[Mux.scala 19:72:@8455.4]
  wire [15:0] _T_5973; // @[Mux.scala 19:72:@8456.4]
  wire [15:0] _T_5974; // @[Mux.scala 19:72:@8457.4]
  wire [15:0] _T_5975; // @[Mux.scala 19:72:@8458.4]
  wire [15:0] _T_5976; // @[Mux.scala 19:72:@8459.4]
  wire [15:0] _T_5977; // @[Mux.scala 19:72:@8460.4]
  wire [15:0] _T_5978; // @[Mux.scala 19:72:@8461.4]
  wire [15:0] _T_5979; // @[Mux.scala 19:72:@8462.4]
  wire [15:0] _T_5980; // @[Mux.scala 19:72:@8463.4]
  wire  _T_6121; // @[LoadQueue.scala 121:105:@8499.4]
  wire  _T_6123; // @[LoadQueue.scala 122:18:@8500.4]
  wire  _T_6125; // @[LoadQueue.scala 122:36:@8501.4]
  wire  _T_6126; // @[LoadQueue.scala 122:27:@8502.4]
  wire  _T_6128; // @[LoadQueue.scala 122:52:@8503.4]
  wire  _T_6130; // @[LoadQueue.scala 122:85:@8504.4]
  wire  _T_6132; // @[LoadQueue.scala 122:103:@8505.4]
  wire  _T_6133; // @[LoadQueue.scala 122:94:@8506.4]
  wire  _T_6135; // @[LoadQueue.scala 122:70:@8507.4]
  wire  _T_6136; // @[LoadQueue.scala 122:67:@8508.4]
  wire  validEntriesInStoreQ_0; // @[LoadQueue.scala 121:91:@8509.4]
  wire  _T_6140; // @[LoadQueue.scala 122:18:@8511.4]
  wire  _T_6142; // @[LoadQueue.scala 122:36:@8512.4]
  wire  _T_6143; // @[LoadQueue.scala 122:27:@8513.4]
  wire  _T_6147; // @[LoadQueue.scala 122:85:@8515.4]
  wire  _T_6149; // @[LoadQueue.scala 122:103:@8516.4]
  wire  _T_6150; // @[LoadQueue.scala 122:94:@8517.4]
  wire  _T_6152; // @[LoadQueue.scala 122:70:@8518.4]
  wire  _T_6153; // @[LoadQueue.scala 122:67:@8519.4]
  wire  validEntriesInStoreQ_1; // @[LoadQueue.scala 121:91:@8520.4]
  wire  _T_6157; // @[LoadQueue.scala 122:18:@8522.4]
  wire  _T_6159; // @[LoadQueue.scala 122:36:@8523.4]
  wire  _T_6160; // @[LoadQueue.scala 122:27:@8524.4]
  wire  _T_6164; // @[LoadQueue.scala 122:85:@8526.4]
  wire  _T_6166; // @[LoadQueue.scala 122:103:@8527.4]
  wire  _T_6167; // @[LoadQueue.scala 122:94:@8528.4]
  wire  _T_6169; // @[LoadQueue.scala 122:70:@8529.4]
  wire  _T_6170; // @[LoadQueue.scala 122:67:@8530.4]
  wire  validEntriesInStoreQ_2; // @[LoadQueue.scala 121:91:@8531.4]
  wire  _T_6174; // @[LoadQueue.scala 122:18:@8533.4]
  wire  _T_6176; // @[LoadQueue.scala 122:36:@8534.4]
  wire  _T_6177; // @[LoadQueue.scala 122:27:@8535.4]
  wire  _T_6181; // @[LoadQueue.scala 122:85:@8537.4]
  wire  _T_6183; // @[LoadQueue.scala 122:103:@8538.4]
  wire  _T_6184; // @[LoadQueue.scala 122:94:@8539.4]
  wire  _T_6186; // @[LoadQueue.scala 122:70:@8540.4]
  wire  _T_6187; // @[LoadQueue.scala 122:67:@8541.4]
  wire  validEntriesInStoreQ_3; // @[LoadQueue.scala 121:91:@8542.4]
  wire  _T_6191; // @[LoadQueue.scala 122:18:@8544.4]
  wire  _T_6193; // @[LoadQueue.scala 122:36:@8545.4]
  wire  _T_6194; // @[LoadQueue.scala 122:27:@8546.4]
  wire  _T_6198; // @[LoadQueue.scala 122:85:@8548.4]
  wire  _T_6200; // @[LoadQueue.scala 122:103:@8549.4]
  wire  _T_6201; // @[LoadQueue.scala 122:94:@8550.4]
  wire  _T_6203; // @[LoadQueue.scala 122:70:@8551.4]
  wire  _T_6204; // @[LoadQueue.scala 122:67:@8552.4]
  wire  validEntriesInStoreQ_4; // @[LoadQueue.scala 121:91:@8553.4]
  wire  _T_6208; // @[LoadQueue.scala 122:18:@8555.4]
  wire  _T_6210; // @[LoadQueue.scala 122:36:@8556.4]
  wire  _T_6211; // @[LoadQueue.scala 122:27:@8557.4]
  wire  _T_6215; // @[LoadQueue.scala 122:85:@8559.4]
  wire  _T_6217; // @[LoadQueue.scala 122:103:@8560.4]
  wire  _T_6218; // @[LoadQueue.scala 122:94:@8561.4]
  wire  _T_6220; // @[LoadQueue.scala 122:70:@8562.4]
  wire  _T_6221; // @[LoadQueue.scala 122:67:@8563.4]
  wire  validEntriesInStoreQ_5; // @[LoadQueue.scala 121:91:@8564.4]
  wire  _T_6225; // @[LoadQueue.scala 122:18:@8566.4]
  wire  _T_6227; // @[LoadQueue.scala 122:36:@8567.4]
  wire  _T_6228; // @[LoadQueue.scala 122:27:@8568.4]
  wire  _T_6232; // @[LoadQueue.scala 122:85:@8570.4]
  wire  _T_6234; // @[LoadQueue.scala 122:103:@8571.4]
  wire  _T_6235; // @[LoadQueue.scala 122:94:@8572.4]
  wire  _T_6237; // @[LoadQueue.scala 122:70:@8573.4]
  wire  _T_6238; // @[LoadQueue.scala 122:67:@8574.4]
  wire  validEntriesInStoreQ_6; // @[LoadQueue.scala 121:91:@8575.4]
  wire  _T_6242; // @[LoadQueue.scala 122:18:@8577.4]
  wire  _T_6244; // @[LoadQueue.scala 122:36:@8578.4]
  wire  _T_6245; // @[LoadQueue.scala 122:27:@8579.4]
  wire  _T_6249; // @[LoadQueue.scala 122:85:@8581.4]
  wire  _T_6251; // @[LoadQueue.scala 122:103:@8582.4]
  wire  _T_6252; // @[LoadQueue.scala 122:94:@8583.4]
  wire  _T_6254; // @[LoadQueue.scala 122:70:@8584.4]
  wire  _T_6255; // @[LoadQueue.scala 122:67:@8585.4]
  wire  validEntriesInStoreQ_7; // @[LoadQueue.scala 121:91:@8586.4]
  wire  _T_6259; // @[LoadQueue.scala 122:18:@8588.4]
  wire  _T_6261; // @[LoadQueue.scala 122:36:@8589.4]
  wire  _T_6262; // @[LoadQueue.scala 122:27:@8590.4]
  wire  _T_6266; // @[LoadQueue.scala 122:85:@8592.4]
  wire  _T_6268; // @[LoadQueue.scala 122:103:@8593.4]
  wire  _T_6269; // @[LoadQueue.scala 122:94:@8594.4]
  wire  _T_6271; // @[LoadQueue.scala 122:70:@8595.4]
  wire  _T_6272; // @[LoadQueue.scala 122:67:@8596.4]
  wire  validEntriesInStoreQ_8; // @[LoadQueue.scala 121:91:@8597.4]
  wire  _T_6276; // @[LoadQueue.scala 122:18:@8599.4]
  wire  _T_6278; // @[LoadQueue.scala 122:36:@8600.4]
  wire  _T_6279; // @[LoadQueue.scala 122:27:@8601.4]
  wire  _T_6283; // @[LoadQueue.scala 122:85:@8603.4]
  wire  _T_6285; // @[LoadQueue.scala 122:103:@8604.4]
  wire  _T_6286; // @[LoadQueue.scala 122:94:@8605.4]
  wire  _T_6288; // @[LoadQueue.scala 122:70:@8606.4]
  wire  _T_6289; // @[LoadQueue.scala 122:67:@8607.4]
  wire  validEntriesInStoreQ_9; // @[LoadQueue.scala 121:91:@8608.4]
  wire  _T_6293; // @[LoadQueue.scala 122:18:@8610.4]
  wire  _T_6295; // @[LoadQueue.scala 122:36:@8611.4]
  wire  _T_6296; // @[LoadQueue.scala 122:27:@8612.4]
  wire  _T_6300; // @[LoadQueue.scala 122:85:@8614.4]
  wire  _T_6302; // @[LoadQueue.scala 122:103:@8615.4]
  wire  _T_6303; // @[LoadQueue.scala 122:94:@8616.4]
  wire  _T_6305; // @[LoadQueue.scala 122:70:@8617.4]
  wire  _T_6306; // @[LoadQueue.scala 122:67:@8618.4]
  wire  validEntriesInStoreQ_10; // @[LoadQueue.scala 121:91:@8619.4]
  wire  _T_6310; // @[LoadQueue.scala 122:18:@8621.4]
  wire  _T_6312; // @[LoadQueue.scala 122:36:@8622.4]
  wire  _T_6313; // @[LoadQueue.scala 122:27:@8623.4]
  wire  _T_6317; // @[LoadQueue.scala 122:85:@8625.4]
  wire  _T_6319; // @[LoadQueue.scala 122:103:@8626.4]
  wire  _T_6320; // @[LoadQueue.scala 122:94:@8627.4]
  wire  _T_6322; // @[LoadQueue.scala 122:70:@8628.4]
  wire  _T_6323; // @[LoadQueue.scala 122:67:@8629.4]
  wire  validEntriesInStoreQ_11; // @[LoadQueue.scala 121:91:@8630.4]
  wire  _T_6327; // @[LoadQueue.scala 122:18:@8632.4]
  wire  _T_6329; // @[LoadQueue.scala 122:36:@8633.4]
  wire  _T_6330; // @[LoadQueue.scala 122:27:@8634.4]
  wire  _T_6334; // @[LoadQueue.scala 122:85:@8636.4]
  wire  _T_6336; // @[LoadQueue.scala 122:103:@8637.4]
  wire  _T_6337; // @[LoadQueue.scala 122:94:@8638.4]
  wire  _T_6339; // @[LoadQueue.scala 122:70:@8639.4]
  wire  _T_6340; // @[LoadQueue.scala 122:67:@8640.4]
  wire  validEntriesInStoreQ_12; // @[LoadQueue.scala 121:91:@8641.4]
  wire  _T_6344; // @[LoadQueue.scala 122:18:@8643.4]
  wire  _T_6346; // @[LoadQueue.scala 122:36:@8644.4]
  wire  _T_6347; // @[LoadQueue.scala 122:27:@8645.4]
  wire  _T_6351; // @[LoadQueue.scala 122:85:@8647.4]
  wire  _T_6353; // @[LoadQueue.scala 122:103:@8648.4]
  wire  _T_6354; // @[LoadQueue.scala 122:94:@8649.4]
  wire  _T_6356; // @[LoadQueue.scala 122:70:@8650.4]
  wire  _T_6357; // @[LoadQueue.scala 122:67:@8651.4]
  wire  validEntriesInStoreQ_13; // @[LoadQueue.scala 121:91:@8652.4]
  wire  _T_6361; // @[LoadQueue.scala 122:18:@8654.4]
  wire  _T_6363; // @[LoadQueue.scala 122:36:@8655.4]
  wire  _T_6364; // @[LoadQueue.scala 122:27:@8656.4]
  wire  _T_6368; // @[LoadQueue.scala 122:85:@8658.4]
  wire  _T_6370; // @[LoadQueue.scala 122:103:@8659.4]
  wire  _T_6371; // @[LoadQueue.scala 122:94:@8660.4]
  wire  _T_6373; // @[LoadQueue.scala 122:70:@8661.4]
  wire  _T_6374; // @[LoadQueue.scala 122:67:@8662.4]
  wire  validEntriesInStoreQ_14; // @[LoadQueue.scala 121:91:@8663.4]
  wire  validEntriesInStoreQ_15; // @[LoadQueue.scala 121:91:@8674.4]
  wire  storesToCheck_0_0; // @[LoadQueue.scala 131:10:@8701.4]
  wire  _T_7662; // @[LoadQueue.scala 131:81:@8704.4]
  wire  _T_7663; // @[LoadQueue.scala 131:72:@8705.4]
  wire  _T_7665; // @[LoadQueue.scala 132:33:@8706.4]
  wire  _T_7668; // @[LoadQueue.scala 132:41:@8708.4]
  wire  _T_7670; // @[LoadQueue.scala 132:9:@8709.4]
  wire  storesToCheck_0_1; // @[LoadQueue.scala 131:10:@8710.4]
  wire  _T_7676; // @[LoadQueue.scala 131:81:@8713.4]
  wire  _T_7677; // @[LoadQueue.scala 131:72:@8714.4]
  wire  _T_7679; // @[LoadQueue.scala 132:33:@8715.4]
  wire  _T_7682; // @[LoadQueue.scala 132:41:@8717.4]
  wire  _T_7684; // @[LoadQueue.scala 132:9:@8718.4]
  wire  storesToCheck_0_2; // @[LoadQueue.scala 131:10:@8719.4]
  wire  _T_7690; // @[LoadQueue.scala 131:81:@8722.4]
  wire  _T_7691; // @[LoadQueue.scala 131:72:@8723.4]
  wire  _T_7693; // @[LoadQueue.scala 132:33:@8724.4]
  wire  _T_7696; // @[LoadQueue.scala 132:41:@8726.4]
  wire  _T_7698; // @[LoadQueue.scala 132:9:@8727.4]
  wire  storesToCheck_0_3; // @[LoadQueue.scala 131:10:@8728.4]
  wire  _T_7704; // @[LoadQueue.scala 131:81:@8731.4]
  wire  _T_7705; // @[LoadQueue.scala 131:72:@8732.4]
  wire  _T_7707; // @[LoadQueue.scala 132:33:@8733.4]
  wire  _T_7710; // @[LoadQueue.scala 132:41:@8735.4]
  wire  _T_7712; // @[LoadQueue.scala 132:9:@8736.4]
  wire  storesToCheck_0_4; // @[LoadQueue.scala 131:10:@8737.4]
  wire  _T_7718; // @[LoadQueue.scala 131:81:@8740.4]
  wire  _T_7719; // @[LoadQueue.scala 131:72:@8741.4]
  wire  _T_7721; // @[LoadQueue.scala 132:33:@8742.4]
  wire  _T_7724; // @[LoadQueue.scala 132:41:@8744.4]
  wire  _T_7726; // @[LoadQueue.scala 132:9:@8745.4]
  wire  storesToCheck_0_5; // @[LoadQueue.scala 131:10:@8746.4]
  wire  _T_7732; // @[LoadQueue.scala 131:81:@8749.4]
  wire  _T_7733; // @[LoadQueue.scala 131:72:@8750.4]
  wire  _T_7735; // @[LoadQueue.scala 132:33:@8751.4]
  wire  _T_7738; // @[LoadQueue.scala 132:41:@8753.4]
  wire  _T_7740; // @[LoadQueue.scala 132:9:@8754.4]
  wire  storesToCheck_0_6; // @[LoadQueue.scala 131:10:@8755.4]
  wire  _T_7746; // @[LoadQueue.scala 131:81:@8758.4]
  wire  _T_7747; // @[LoadQueue.scala 131:72:@8759.4]
  wire  _T_7749; // @[LoadQueue.scala 132:33:@8760.4]
  wire  _T_7752; // @[LoadQueue.scala 132:41:@8762.4]
  wire  _T_7754; // @[LoadQueue.scala 132:9:@8763.4]
  wire  storesToCheck_0_7; // @[LoadQueue.scala 131:10:@8764.4]
  wire  _T_7760; // @[LoadQueue.scala 131:81:@8767.4]
  wire  _T_7761; // @[LoadQueue.scala 131:72:@8768.4]
  wire  _T_7763; // @[LoadQueue.scala 132:33:@8769.4]
  wire  _T_7766; // @[LoadQueue.scala 132:41:@8771.4]
  wire  _T_7768; // @[LoadQueue.scala 132:9:@8772.4]
  wire  storesToCheck_0_8; // @[LoadQueue.scala 131:10:@8773.4]
  wire  _T_7774; // @[LoadQueue.scala 131:81:@8776.4]
  wire  _T_7775; // @[LoadQueue.scala 131:72:@8777.4]
  wire  _T_7777; // @[LoadQueue.scala 132:33:@8778.4]
  wire  _T_7780; // @[LoadQueue.scala 132:41:@8780.4]
  wire  _T_7782; // @[LoadQueue.scala 132:9:@8781.4]
  wire  storesToCheck_0_9; // @[LoadQueue.scala 131:10:@8782.4]
  wire  _T_7788; // @[LoadQueue.scala 131:81:@8785.4]
  wire  _T_7789; // @[LoadQueue.scala 131:72:@8786.4]
  wire  _T_7791; // @[LoadQueue.scala 132:33:@8787.4]
  wire  _T_7794; // @[LoadQueue.scala 132:41:@8789.4]
  wire  _T_7796; // @[LoadQueue.scala 132:9:@8790.4]
  wire  storesToCheck_0_10; // @[LoadQueue.scala 131:10:@8791.4]
  wire  _T_7802; // @[LoadQueue.scala 131:81:@8794.4]
  wire  _T_7803; // @[LoadQueue.scala 131:72:@8795.4]
  wire  _T_7805; // @[LoadQueue.scala 132:33:@8796.4]
  wire  _T_7808; // @[LoadQueue.scala 132:41:@8798.4]
  wire  _T_7810; // @[LoadQueue.scala 132:9:@8799.4]
  wire  storesToCheck_0_11; // @[LoadQueue.scala 131:10:@8800.4]
  wire  _T_7816; // @[LoadQueue.scala 131:81:@8803.4]
  wire  _T_7817; // @[LoadQueue.scala 131:72:@8804.4]
  wire  _T_7819; // @[LoadQueue.scala 132:33:@8805.4]
  wire  _T_7822; // @[LoadQueue.scala 132:41:@8807.4]
  wire  _T_7824; // @[LoadQueue.scala 132:9:@8808.4]
  wire  storesToCheck_0_12; // @[LoadQueue.scala 131:10:@8809.4]
  wire  _T_7830; // @[LoadQueue.scala 131:81:@8812.4]
  wire  _T_7831; // @[LoadQueue.scala 131:72:@8813.4]
  wire  _T_7833; // @[LoadQueue.scala 132:33:@8814.4]
  wire  _T_7836; // @[LoadQueue.scala 132:41:@8816.4]
  wire  _T_7838; // @[LoadQueue.scala 132:9:@8817.4]
  wire  storesToCheck_0_13; // @[LoadQueue.scala 131:10:@8818.4]
  wire  _T_7844; // @[LoadQueue.scala 131:81:@8821.4]
  wire  _T_7845; // @[LoadQueue.scala 131:72:@8822.4]
  wire  _T_7847; // @[LoadQueue.scala 132:33:@8823.4]
  wire  _T_7850; // @[LoadQueue.scala 132:41:@8825.4]
  wire  _T_7852; // @[LoadQueue.scala 132:9:@8826.4]
  wire  storesToCheck_0_14; // @[LoadQueue.scala 131:10:@8827.4]
  wire  _T_7858; // @[LoadQueue.scala 131:81:@8830.4]
  wire  storesToCheck_0_15; // @[LoadQueue.scala 131:10:@8836.4]
  wire  storesToCheck_1_0; // @[LoadQueue.scala 131:10:@8878.4]
  wire  _T_7908; // @[LoadQueue.scala 131:81:@8881.4]
  wire  _T_7909; // @[LoadQueue.scala 131:72:@8882.4]
  wire  _T_7911; // @[LoadQueue.scala 132:33:@8883.4]
  wire  _T_7914; // @[LoadQueue.scala 132:41:@8885.4]
  wire  _T_7916; // @[LoadQueue.scala 132:9:@8886.4]
  wire  storesToCheck_1_1; // @[LoadQueue.scala 131:10:@8887.4]
  wire  _T_7922; // @[LoadQueue.scala 131:81:@8890.4]
  wire  _T_7923; // @[LoadQueue.scala 131:72:@8891.4]
  wire  _T_7925; // @[LoadQueue.scala 132:33:@8892.4]
  wire  _T_7928; // @[LoadQueue.scala 132:41:@8894.4]
  wire  _T_7930; // @[LoadQueue.scala 132:9:@8895.4]
  wire  storesToCheck_1_2; // @[LoadQueue.scala 131:10:@8896.4]
  wire  _T_7936; // @[LoadQueue.scala 131:81:@8899.4]
  wire  _T_7937; // @[LoadQueue.scala 131:72:@8900.4]
  wire  _T_7939; // @[LoadQueue.scala 132:33:@8901.4]
  wire  _T_7942; // @[LoadQueue.scala 132:41:@8903.4]
  wire  _T_7944; // @[LoadQueue.scala 132:9:@8904.4]
  wire  storesToCheck_1_3; // @[LoadQueue.scala 131:10:@8905.4]
  wire  _T_7950; // @[LoadQueue.scala 131:81:@8908.4]
  wire  _T_7951; // @[LoadQueue.scala 131:72:@8909.4]
  wire  _T_7953; // @[LoadQueue.scala 132:33:@8910.4]
  wire  _T_7956; // @[LoadQueue.scala 132:41:@8912.4]
  wire  _T_7958; // @[LoadQueue.scala 132:9:@8913.4]
  wire  storesToCheck_1_4; // @[LoadQueue.scala 131:10:@8914.4]
  wire  _T_7964; // @[LoadQueue.scala 131:81:@8917.4]
  wire  _T_7965; // @[LoadQueue.scala 131:72:@8918.4]
  wire  _T_7967; // @[LoadQueue.scala 132:33:@8919.4]
  wire  _T_7970; // @[LoadQueue.scala 132:41:@8921.4]
  wire  _T_7972; // @[LoadQueue.scala 132:9:@8922.4]
  wire  storesToCheck_1_5; // @[LoadQueue.scala 131:10:@8923.4]
  wire  _T_7978; // @[LoadQueue.scala 131:81:@8926.4]
  wire  _T_7979; // @[LoadQueue.scala 131:72:@8927.4]
  wire  _T_7981; // @[LoadQueue.scala 132:33:@8928.4]
  wire  _T_7984; // @[LoadQueue.scala 132:41:@8930.4]
  wire  _T_7986; // @[LoadQueue.scala 132:9:@8931.4]
  wire  storesToCheck_1_6; // @[LoadQueue.scala 131:10:@8932.4]
  wire  _T_7992; // @[LoadQueue.scala 131:81:@8935.4]
  wire  _T_7993; // @[LoadQueue.scala 131:72:@8936.4]
  wire  _T_7995; // @[LoadQueue.scala 132:33:@8937.4]
  wire  _T_7998; // @[LoadQueue.scala 132:41:@8939.4]
  wire  _T_8000; // @[LoadQueue.scala 132:9:@8940.4]
  wire  storesToCheck_1_7; // @[LoadQueue.scala 131:10:@8941.4]
  wire  _T_8006; // @[LoadQueue.scala 131:81:@8944.4]
  wire  _T_8007; // @[LoadQueue.scala 131:72:@8945.4]
  wire  _T_8009; // @[LoadQueue.scala 132:33:@8946.4]
  wire  _T_8012; // @[LoadQueue.scala 132:41:@8948.4]
  wire  _T_8014; // @[LoadQueue.scala 132:9:@8949.4]
  wire  storesToCheck_1_8; // @[LoadQueue.scala 131:10:@8950.4]
  wire  _T_8020; // @[LoadQueue.scala 131:81:@8953.4]
  wire  _T_8021; // @[LoadQueue.scala 131:72:@8954.4]
  wire  _T_8023; // @[LoadQueue.scala 132:33:@8955.4]
  wire  _T_8026; // @[LoadQueue.scala 132:41:@8957.4]
  wire  _T_8028; // @[LoadQueue.scala 132:9:@8958.4]
  wire  storesToCheck_1_9; // @[LoadQueue.scala 131:10:@8959.4]
  wire  _T_8034; // @[LoadQueue.scala 131:81:@8962.4]
  wire  _T_8035; // @[LoadQueue.scala 131:72:@8963.4]
  wire  _T_8037; // @[LoadQueue.scala 132:33:@8964.4]
  wire  _T_8040; // @[LoadQueue.scala 132:41:@8966.4]
  wire  _T_8042; // @[LoadQueue.scala 132:9:@8967.4]
  wire  storesToCheck_1_10; // @[LoadQueue.scala 131:10:@8968.4]
  wire  _T_8048; // @[LoadQueue.scala 131:81:@8971.4]
  wire  _T_8049; // @[LoadQueue.scala 131:72:@8972.4]
  wire  _T_8051; // @[LoadQueue.scala 132:33:@8973.4]
  wire  _T_8054; // @[LoadQueue.scala 132:41:@8975.4]
  wire  _T_8056; // @[LoadQueue.scala 132:9:@8976.4]
  wire  storesToCheck_1_11; // @[LoadQueue.scala 131:10:@8977.4]
  wire  _T_8062; // @[LoadQueue.scala 131:81:@8980.4]
  wire  _T_8063; // @[LoadQueue.scala 131:72:@8981.4]
  wire  _T_8065; // @[LoadQueue.scala 132:33:@8982.4]
  wire  _T_8068; // @[LoadQueue.scala 132:41:@8984.4]
  wire  _T_8070; // @[LoadQueue.scala 132:9:@8985.4]
  wire  storesToCheck_1_12; // @[LoadQueue.scala 131:10:@8986.4]
  wire  _T_8076; // @[LoadQueue.scala 131:81:@8989.4]
  wire  _T_8077; // @[LoadQueue.scala 131:72:@8990.4]
  wire  _T_8079; // @[LoadQueue.scala 132:33:@8991.4]
  wire  _T_8082; // @[LoadQueue.scala 132:41:@8993.4]
  wire  _T_8084; // @[LoadQueue.scala 132:9:@8994.4]
  wire  storesToCheck_1_13; // @[LoadQueue.scala 131:10:@8995.4]
  wire  _T_8090; // @[LoadQueue.scala 131:81:@8998.4]
  wire  _T_8091; // @[LoadQueue.scala 131:72:@8999.4]
  wire  _T_8093; // @[LoadQueue.scala 132:33:@9000.4]
  wire  _T_8096; // @[LoadQueue.scala 132:41:@9002.4]
  wire  _T_8098; // @[LoadQueue.scala 132:9:@9003.4]
  wire  storesToCheck_1_14; // @[LoadQueue.scala 131:10:@9004.4]
  wire  _T_8104; // @[LoadQueue.scala 131:81:@9007.4]
  wire  storesToCheck_1_15; // @[LoadQueue.scala 131:10:@9013.4]
  wire  storesToCheck_2_0; // @[LoadQueue.scala 131:10:@9055.4]
  wire  _T_8154; // @[LoadQueue.scala 131:81:@9058.4]
  wire  _T_8155; // @[LoadQueue.scala 131:72:@9059.4]
  wire  _T_8157; // @[LoadQueue.scala 132:33:@9060.4]
  wire  _T_8160; // @[LoadQueue.scala 132:41:@9062.4]
  wire  _T_8162; // @[LoadQueue.scala 132:9:@9063.4]
  wire  storesToCheck_2_1; // @[LoadQueue.scala 131:10:@9064.4]
  wire  _T_8168; // @[LoadQueue.scala 131:81:@9067.4]
  wire  _T_8169; // @[LoadQueue.scala 131:72:@9068.4]
  wire  _T_8171; // @[LoadQueue.scala 132:33:@9069.4]
  wire  _T_8174; // @[LoadQueue.scala 132:41:@9071.4]
  wire  _T_8176; // @[LoadQueue.scala 132:9:@9072.4]
  wire  storesToCheck_2_2; // @[LoadQueue.scala 131:10:@9073.4]
  wire  _T_8182; // @[LoadQueue.scala 131:81:@9076.4]
  wire  _T_8183; // @[LoadQueue.scala 131:72:@9077.4]
  wire  _T_8185; // @[LoadQueue.scala 132:33:@9078.4]
  wire  _T_8188; // @[LoadQueue.scala 132:41:@9080.4]
  wire  _T_8190; // @[LoadQueue.scala 132:9:@9081.4]
  wire  storesToCheck_2_3; // @[LoadQueue.scala 131:10:@9082.4]
  wire  _T_8196; // @[LoadQueue.scala 131:81:@9085.4]
  wire  _T_8197; // @[LoadQueue.scala 131:72:@9086.4]
  wire  _T_8199; // @[LoadQueue.scala 132:33:@9087.4]
  wire  _T_8202; // @[LoadQueue.scala 132:41:@9089.4]
  wire  _T_8204; // @[LoadQueue.scala 132:9:@9090.4]
  wire  storesToCheck_2_4; // @[LoadQueue.scala 131:10:@9091.4]
  wire  _T_8210; // @[LoadQueue.scala 131:81:@9094.4]
  wire  _T_8211; // @[LoadQueue.scala 131:72:@9095.4]
  wire  _T_8213; // @[LoadQueue.scala 132:33:@9096.4]
  wire  _T_8216; // @[LoadQueue.scala 132:41:@9098.4]
  wire  _T_8218; // @[LoadQueue.scala 132:9:@9099.4]
  wire  storesToCheck_2_5; // @[LoadQueue.scala 131:10:@9100.4]
  wire  _T_8224; // @[LoadQueue.scala 131:81:@9103.4]
  wire  _T_8225; // @[LoadQueue.scala 131:72:@9104.4]
  wire  _T_8227; // @[LoadQueue.scala 132:33:@9105.4]
  wire  _T_8230; // @[LoadQueue.scala 132:41:@9107.4]
  wire  _T_8232; // @[LoadQueue.scala 132:9:@9108.4]
  wire  storesToCheck_2_6; // @[LoadQueue.scala 131:10:@9109.4]
  wire  _T_8238; // @[LoadQueue.scala 131:81:@9112.4]
  wire  _T_8239; // @[LoadQueue.scala 131:72:@9113.4]
  wire  _T_8241; // @[LoadQueue.scala 132:33:@9114.4]
  wire  _T_8244; // @[LoadQueue.scala 132:41:@9116.4]
  wire  _T_8246; // @[LoadQueue.scala 132:9:@9117.4]
  wire  storesToCheck_2_7; // @[LoadQueue.scala 131:10:@9118.4]
  wire  _T_8252; // @[LoadQueue.scala 131:81:@9121.4]
  wire  _T_8253; // @[LoadQueue.scala 131:72:@9122.4]
  wire  _T_8255; // @[LoadQueue.scala 132:33:@9123.4]
  wire  _T_8258; // @[LoadQueue.scala 132:41:@9125.4]
  wire  _T_8260; // @[LoadQueue.scala 132:9:@9126.4]
  wire  storesToCheck_2_8; // @[LoadQueue.scala 131:10:@9127.4]
  wire  _T_8266; // @[LoadQueue.scala 131:81:@9130.4]
  wire  _T_8267; // @[LoadQueue.scala 131:72:@9131.4]
  wire  _T_8269; // @[LoadQueue.scala 132:33:@9132.4]
  wire  _T_8272; // @[LoadQueue.scala 132:41:@9134.4]
  wire  _T_8274; // @[LoadQueue.scala 132:9:@9135.4]
  wire  storesToCheck_2_9; // @[LoadQueue.scala 131:10:@9136.4]
  wire  _T_8280; // @[LoadQueue.scala 131:81:@9139.4]
  wire  _T_8281; // @[LoadQueue.scala 131:72:@9140.4]
  wire  _T_8283; // @[LoadQueue.scala 132:33:@9141.4]
  wire  _T_8286; // @[LoadQueue.scala 132:41:@9143.4]
  wire  _T_8288; // @[LoadQueue.scala 132:9:@9144.4]
  wire  storesToCheck_2_10; // @[LoadQueue.scala 131:10:@9145.4]
  wire  _T_8294; // @[LoadQueue.scala 131:81:@9148.4]
  wire  _T_8295; // @[LoadQueue.scala 131:72:@9149.4]
  wire  _T_8297; // @[LoadQueue.scala 132:33:@9150.4]
  wire  _T_8300; // @[LoadQueue.scala 132:41:@9152.4]
  wire  _T_8302; // @[LoadQueue.scala 132:9:@9153.4]
  wire  storesToCheck_2_11; // @[LoadQueue.scala 131:10:@9154.4]
  wire  _T_8308; // @[LoadQueue.scala 131:81:@9157.4]
  wire  _T_8309; // @[LoadQueue.scala 131:72:@9158.4]
  wire  _T_8311; // @[LoadQueue.scala 132:33:@9159.4]
  wire  _T_8314; // @[LoadQueue.scala 132:41:@9161.4]
  wire  _T_8316; // @[LoadQueue.scala 132:9:@9162.4]
  wire  storesToCheck_2_12; // @[LoadQueue.scala 131:10:@9163.4]
  wire  _T_8322; // @[LoadQueue.scala 131:81:@9166.4]
  wire  _T_8323; // @[LoadQueue.scala 131:72:@9167.4]
  wire  _T_8325; // @[LoadQueue.scala 132:33:@9168.4]
  wire  _T_8328; // @[LoadQueue.scala 132:41:@9170.4]
  wire  _T_8330; // @[LoadQueue.scala 132:9:@9171.4]
  wire  storesToCheck_2_13; // @[LoadQueue.scala 131:10:@9172.4]
  wire  _T_8336; // @[LoadQueue.scala 131:81:@9175.4]
  wire  _T_8337; // @[LoadQueue.scala 131:72:@9176.4]
  wire  _T_8339; // @[LoadQueue.scala 132:33:@9177.4]
  wire  _T_8342; // @[LoadQueue.scala 132:41:@9179.4]
  wire  _T_8344; // @[LoadQueue.scala 132:9:@9180.4]
  wire  storesToCheck_2_14; // @[LoadQueue.scala 131:10:@9181.4]
  wire  _T_8350; // @[LoadQueue.scala 131:81:@9184.4]
  wire  storesToCheck_2_15; // @[LoadQueue.scala 131:10:@9190.4]
  wire  storesToCheck_3_0; // @[LoadQueue.scala 131:10:@9232.4]
  wire  _T_8400; // @[LoadQueue.scala 131:81:@9235.4]
  wire  _T_8401; // @[LoadQueue.scala 131:72:@9236.4]
  wire  _T_8403; // @[LoadQueue.scala 132:33:@9237.4]
  wire  _T_8406; // @[LoadQueue.scala 132:41:@9239.4]
  wire  _T_8408; // @[LoadQueue.scala 132:9:@9240.4]
  wire  storesToCheck_3_1; // @[LoadQueue.scala 131:10:@9241.4]
  wire  _T_8414; // @[LoadQueue.scala 131:81:@9244.4]
  wire  _T_8415; // @[LoadQueue.scala 131:72:@9245.4]
  wire  _T_8417; // @[LoadQueue.scala 132:33:@9246.4]
  wire  _T_8420; // @[LoadQueue.scala 132:41:@9248.4]
  wire  _T_8422; // @[LoadQueue.scala 132:9:@9249.4]
  wire  storesToCheck_3_2; // @[LoadQueue.scala 131:10:@9250.4]
  wire  _T_8428; // @[LoadQueue.scala 131:81:@9253.4]
  wire  _T_8429; // @[LoadQueue.scala 131:72:@9254.4]
  wire  _T_8431; // @[LoadQueue.scala 132:33:@9255.4]
  wire  _T_8434; // @[LoadQueue.scala 132:41:@9257.4]
  wire  _T_8436; // @[LoadQueue.scala 132:9:@9258.4]
  wire  storesToCheck_3_3; // @[LoadQueue.scala 131:10:@9259.4]
  wire  _T_8442; // @[LoadQueue.scala 131:81:@9262.4]
  wire  _T_8443; // @[LoadQueue.scala 131:72:@9263.4]
  wire  _T_8445; // @[LoadQueue.scala 132:33:@9264.4]
  wire  _T_8448; // @[LoadQueue.scala 132:41:@9266.4]
  wire  _T_8450; // @[LoadQueue.scala 132:9:@9267.4]
  wire  storesToCheck_3_4; // @[LoadQueue.scala 131:10:@9268.4]
  wire  _T_8456; // @[LoadQueue.scala 131:81:@9271.4]
  wire  _T_8457; // @[LoadQueue.scala 131:72:@9272.4]
  wire  _T_8459; // @[LoadQueue.scala 132:33:@9273.4]
  wire  _T_8462; // @[LoadQueue.scala 132:41:@9275.4]
  wire  _T_8464; // @[LoadQueue.scala 132:9:@9276.4]
  wire  storesToCheck_3_5; // @[LoadQueue.scala 131:10:@9277.4]
  wire  _T_8470; // @[LoadQueue.scala 131:81:@9280.4]
  wire  _T_8471; // @[LoadQueue.scala 131:72:@9281.4]
  wire  _T_8473; // @[LoadQueue.scala 132:33:@9282.4]
  wire  _T_8476; // @[LoadQueue.scala 132:41:@9284.4]
  wire  _T_8478; // @[LoadQueue.scala 132:9:@9285.4]
  wire  storesToCheck_3_6; // @[LoadQueue.scala 131:10:@9286.4]
  wire  _T_8484; // @[LoadQueue.scala 131:81:@9289.4]
  wire  _T_8485; // @[LoadQueue.scala 131:72:@9290.4]
  wire  _T_8487; // @[LoadQueue.scala 132:33:@9291.4]
  wire  _T_8490; // @[LoadQueue.scala 132:41:@9293.4]
  wire  _T_8492; // @[LoadQueue.scala 132:9:@9294.4]
  wire  storesToCheck_3_7; // @[LoadQueue.scala 131:10:@9295.4]
  wire  _T_8498; // @[LoadQueue.scala 131:81:@9298.4]
  wire  _T_8499; // @[LoadQueue.scala 131:72:@9299.4]
  wire  _T_8501; // @[LoadQueue.scala 132:33:@9300.4]
  wire  _T_8504; // @[LoadQueue.scala 132:41:@9302.4]
  wire  _T_8506; // @[LoadQueue.scala 132:9:@9303.4]
  wire  storesToCheck_3_8; // @[LoadQueue.scala 131:10:@9304.4]
  wire  _T_8512; // @[LoadQueue.scala 131:81:@9307.4]
  wire  _T_8513; // @[LoadQueue.scala 131:72:@9308.4]
  wire  _T_8515; // @[LoadQueue.scala 132:33:@9309.4]
  wire  _T_8518; // @[LoadQueue.scala 132:41:@9311.4]
  wire  _T_8520; // @[LoadQueue.scala 132:9:@9312.4]
  wire  storesToCheck_3_9; // @[LoadQueue.scala 131:10:@9313.4]
  wire  _T_8526; // @[LoadQueue.scala 131:81:@9316.4]
  wire  _T_8527; // @[LoadQueue.scala 131:72:@9317.4]
  wire  _T_8529; // @[LoadQueue.scala 132:33:@9318.4]
  wire  _T_8532; // @[LoadQueue.scala 132:41:@9320.4]
  wire  _T_8534; // @[LoadQueue.scala 132:9:@9321.4]
  wire  storesToCheck_3_10; // @[LoadQueue.scala 131:10:@9322.4]
  wire  _T_8540; // @[LoadQueue.scala 131:81:@9325.4]
  wire  _T_8541; // @[LoadQueue.scala 131:72:@9326.4]
  wire  _T_8543; // @[LoadQueue.scala 132:33:@9327.4]
  wire  _T_8546; // @[LoadQueue.scala 132:41:@9329.4]
  wire  _T_8548; // @[LoadQueue.scala 132:9:@9330.4]
  wire  storesToCheck_3_11; // @[LoadQueue.scala 131:10:@9331.4]
  wire  _T_8554; // @[LoadQueue.scala 131:81:@9334.4]
  wire  _T_8555; // @[LoadQueue.scala 131:72:@9335.4]
  wire  _T_8557; // @[LoadQueue.scala 132:33:@9336.4]
  wire  _T_8560; // @[LoadQueue.scala 132:41:@9338.4]
  wire  _T_8562; // @[LoadQueue.scala 132:9:@9339.4]
  wire  storesToCheck_3_12; // @[LoadQueue.scala 131:10:@9340.4]
  wire  _T_8568; // @[LoadQueue.scala 131:81:@9343.4]
  wire  _T_8569; // @[LoadQueue.scala 131:72:@9344.4]
  wire  _T_8571; // @[LoadQueue.scala 132:33:@9345.4]
  wire  _T_8574; // @[LoadQueue.scala 132:41:@9347.4]
  wire  _T_8576; // @[LoadQueue.scala 132:9:@9348.4]
  wire  storesToCheck_3_13; // @[LoadQueue.scala 131:10:@9349.4]
  wire  _T_8582; // @[LoadQueue.scala 131:81:@9352.4]
  wire  _T_8583; // @[LoadQueue.scala 131:72:@9353.4]
  wire  _T_8585; // @[LoadQueue.scala 132:33:@9354.4]
  wire  _T_8588; // @[LoadQueue.scala 132:41:@9356.4]
  wire  _T_8590; // @[LoadQueue.scala 132:9:@9357.4]
  wire  storesToCheck_3_14; // @[LoadQueue.scala 131:10:@9358.4]
  wire  _T_8596; // @[LoadQueue.scala 131:81:@9361.4]
  wire  storesToCheck_3_15; // @[LoadQueue.scala 131:10:@9367.4]
  wire  storesToCheck_4_0; // @[LoadQueue.scala 131:10:@9409.4]
  wire  _T_8646; // @[LoadQueue.scala 131:81:@9412.4]
  wire  _T_8647; // @[LoadQueue.scala 131:72:@9413.4]
  wire  _T_8649; // @[LoadQueue.scala 132:33:@9414.4]
  wire  _T_8652; // @[LoadQueue.scala 132:41:@9416.4]
  wire  _T_8654; // @[LoadQueue.scala 132:9:@9417.4]
  wire  storesToCheck_4_1; // @[LoadQueue.scala 131:10:@9418.4]
  wire  _T_8660; // @[LoadQueue.scala 131:81:@9421.4]
  wire  _T_8661; // @[LoadQueue.scala 131:72:@9422.4]
  wire  _T_8663; // @[LoadQueue.scala 132:33:@9423.4]
  wire  _T_8666; // @[LoadQueue.scala 132:41:@9425.4]
  wire  _T_8668; // @[LoadQueue.scala 132:9:@9426.4]
  wire  storesToCheck_4_2; // @[LoadQueue.scala 131:10:@9427.4]
  wire  _T_8674; // @[LoadQueue.scala 131:81:@9430.4]
  wire  _T_8675; // @[LoadQueue.scala 131:72:@9431.4]
  wire  _T_8677; // @[LoadQueue.scala 132:33:@9432.4]
  wire  _T_8680; // @[LoadQueue.scala 132:41:@9434.4]
  wire  _T_8682; // @[LoadQueue.scala 132:9:@9435.4]
  wire  storesToCheck_4_3; // @[LoadQueue.scala 131:10:@9436.4]
  wire  _T_8688; // @[LoadQueue.scala 131:81:@9439.4]
  wire  _T_8689; // @[LoadQueue.scala 131:72:@9440.4]
  wire  _T_8691; // @[LoadQueue.scala 132:33:@9441.4]
  wire  _T_8694; // @[LoadQueue.scala 132:41:@9443.4]
  wire  _T_8696; // @[LoadQueue.scala 132:9:@9444.4]
  wire  storesToCheck_4_4; // @[LoadQueue.scala 131:10:@9445.4]
  wire  _T_8702; // @[LoadQueue.scala 131:81:@9448.4]
  wire  _T_8703; // @[LoadQueue.scala 131:72:@9449.4]
  wire  _T_8705; // @[LoadQueue.scala 132:33:@9450.4]
  wire  _T_8708; // @[LoadQueue.scala 132:41:@9452.4]
  wire  _T_8710; // @[LoadQueue.scala 132:9:@9453.4]
  wire  storesToCheck_4_5; // @[LoadQueue.scala 131:10:@9454.4]
  wire  _T_8716; // @[LoadQueue.scala 131:81:@9457.4]
  wire  _T_8717; // @[LoadQueue.scala 131:72:@9458.4]
  wire  _T_8719; // @[LoadQueue.scala 132:33:@9459.4]
  wire  _T_8722; // @[LoadQueue.scala 132:41:@9461.4]
  wire  _T_8724; // @[LoadQueue.scala 132:9:@9462.4]
  wire  storesToCheck_4_6; // @[LoadQueue.scala 131:10:@9463.4]
  wire  _T_8730; // @[LoadQueue.scala 131:81:@9466.4]
  wire  _T_8731; // @[LoadQueue.scala 131:72:@9467.4]
  wire  _T_8733; // @[LoadQueue.scala 132:33:@9468.4]
  wire  _T_8736; // @[LoadQueue.scala 132:41:@9470.4]
  wire  _T_8738; // @[LoadQueue.scala 132:9:@9471.4]
  wire  storesToCheck_4_7; // @[LoadQueue.scala 131:10:@9472.4]
  wire  _T_8744; // @[LoadQueue.scala 131:81:@9475.4]
  wire  _T_8745; // @[LoadQueue.scala 131:72:@9476.4]
  wire  _T_8747; // @[LoadQueue.scala 132:33:@9477.4]
  wire  _T_8750; // @[LoadQueue.scala 132:41:@9479.4]
  wire  _T_8752; // @[LoadQueue.scala 132:9:@9480.4]
  wire  storesToCheck_4_8; // @[LoadQueue.scala 131:10:@9481.4]
  wire  _T_8758; // @[LoadQueue.scala 131:81:@9484.4]
  wire  _T_8759; // @[LoadQueue.scala 131:72:@9485.4]
  wire  _T_8761; // @[LoadQueue.scala 132:33:@9486.4]
  wire  _T_8764; // @[LoadQueue.scala 132:41:@9488.4]
  wire  _T_8766; // @[LoadQueue.scala 132:9:@9489.4]
  wire  storesToCheck_4_9; // @[LoadQueue.scala 131:10:@9490.4]
  wire  _T_8772; // @[LoadQueue.scala 131:81:@9493.4]
  wire  _T_8773; // @[LoadQueue.scala 131:72:@9494.4]
  wire  _T_8775; // @[LoadQueue.scala 132:33:@9495.4]
  wire  _T_8778; // @[LoadQueue.scala 132:41:@9497.4]
  wire  _T_8780; // @[LoadQueue.scala 132:9:@9498.4]
  wire  storesToCheck_4_10; // @[LoadQueue.scala 131:10:@9499.4]
  wire  _T_8786; // @[LoadQueue.scala 131:81:@9502.4]
  wire  _T_8787; // @[LoadQueue.scala 131:72:@9503.4]
  wire  _T_8789; // @[LoadQueue.scala 132:33:@9504.4]
  wire  _T_8792; // @[LoadQueue.scala 132:41:@9506.4]
  wire  _T_8794; // @[LoadQueue.scala 132:9:@9507.4]
  wire  storesToCheck_4_11; // @[LoadQueue.scala 131:10:@9508.4]
  wire  _T_8800; // @[LoadQueue.scala 131:81:@9511.4]
  wire  _T_8801; // @[LoadQueue.scala 131:72:@9512.4]
  wire  _T_8803; // @[LoadQueue.scala 132:33:@9513.4]
  wire  _T_8806; // @[LoadQueue.scala 132:41:@9515.4]
  wire  _T_8808; // @[LoadQueue.scala 132:9:@9516.4]
  wire  storesToCheck_4_12; // @[LoadQueue.scala 131:10:@9517.4]
  wire  _T_8814; // @[LoadQueue.scala 131:81:@9520.4]
  wire  _T_8815; // @[LoadQueue.scala 131:72:@9521.4]
  wire  _T_8817; // @[LoadQueue.scala 132:33:@9522.4]
  wire  _T_8820; // @[LoadQueue.scala 132:41:@9524.4]
  wire  _T_8822; // @[LoadQueue.scala 132:9:@9525.4]
  wire  storesToCheck_4_13; // @[LoadQueue.scala 131:10:@9526.4]
  wire  _T_8828; // @[LoadQueue.scala 131:81:@9529.4]
  wire  _T_8829; // @[LoadQueue.scala 131:72:@9530.4]
  wire  _T_8831; // @[LoadQueue.scala 132:33:@9531.4]
  wire  _T_8834; // @[LoadQueue.scala 132:41:@9533.4]
  wire  _T_8836; // @[LoadQueue.scala 132:9:@9534.4]
  wire  storesToCheck_4_14; // @[LoadQueue.scala 131:10:@9535.4]
  wire  _T_8842; // @[LoadQueue.scala 131:81:@9538.4]
  wire  storesToCheck_4_15; // @[LoadQueue.scala 131:10:@9544.4]
  wire  storesToCheck_5_0; // @[LoadQueue.scala 131:10:@9586.4]
  wire  _T_8892; // @[LoadQueue.scala 131:81:@9589.4]
  wire  _T_8893; // @[LoadQueue.scala 131:72:@9590.4]
  wire  _T_8895; // @[LoadQueue.scala 132:33:@9591.4]
  wire  _T_8898; // @[LoadQueue.scala 132:41:@9593.4]
  wire  _T_8900; // @[LoadQueue.scala 132:9:@9594.4]
  wire  storesToCheck_5_1; // @[LoadQueue.scala 131:10:@9595.4]
  wire  _T_8906; // @[LoadQueue.scala 131:81:@9598.4]
  wire  _T_8907; // @[LoadQueue.scala 131:72:@9599.4]
  wire  _T_8909; // @[LoadQueue.scala 132:33:@9600.4]
  wire  _T_8912; // @[LoadQueue.scala 132:41:@9602.4]
  wire  _T_8914; // @[LoadQueue.scala 132:9:@9603.4]
  wire  storesToCheck_5_2; // @[LoadQueue.scala 131:10:@9604.4]
  wire  _T_8920; // @[LoadQueue.scala 131:81:@9607.4]
  wire  _T_8921; // @[LoadQueue.scala 131:72:@9608.4]
  wire  _T_8923; // @[LoadQueue.scala 132:33:@9609.4]
  wire  _T_8926; // @[LoadQueue.scala 132:41:@9611.4]
  wire  _T_8928; // @[LoadQueue.scala 132:9:@9612.4]
  wire  storesToCheck_5_3; // @[LoadQueue.scala 131:10:@9613.4]
  wire  _T_8934; // @[LoadQueue.scala 131:81:@9616.4]
  wire  _T_8935; // @[LoadQueue.scala 131:72:@9617.4]
  wire  _T_8937; // @[LoadQueue.scala 132:33:@9618.4]
  wire  _T_8940; // @[LoadQueue.scala 132:41:@9620.4]
  wire  _T_8942; // @[LoadQueue.scala 132:9:@9621.4]
  wire  storesToCheck_5_4; // @[LoadQueue.scala 131:10:@9622.4]
  wire  _T_8948; // @[LoadQueue.scala 131:81:@9625.4]
  wire  _T_8949; // @[LoadQueue.scala 131:72:@9626.4]
  wire  _T_8951; // @[LoadQueue.scala 132:33:@9627.4]
  wire  _T_8954; // @[LoadQueue.scala 132:41:@9629.4]
  wire  _T_8956; // @[LoadQueue.scala 132:9:@9630.4]
  wire  storesToCheck_5_5; // @[LoadQueue.scala 131:10:@9631.4]
  wire  _T_8962; // @[LoadQueue.scala 131:81:@9634.4]
  wire  _T_8963; // @[LoadQueue.scala 131:72:@9635.4]
  wire  _T_8965; // @[LoadQueue.scala 132:33:@9636.4]
  wire  _T_8968; // @[LoadQueue.scala 132:41:@9638.4]
  wire  _T_8970; // @[LoadQueue.scala 132:9:@9639.4]
  wire  storesToCheck_5_6; // @[LoadQueue.scala 131:10:@9640.4]
  wire  _T_8976; // @[LoadQueue.scala 131:81:@9643.4]
  wire  _T_8977; // @[LoadQueue.scala 131:72:@9644.4]
  wire  _T_8979; // @[LoadQueue.scala 132:33:@9645.4]
  wire  _T_8982; // @[LoadQueue.scala 132:41:@9647.4]
  wire  _T_8984; // @[LoadQueue.scala 132:9:@9648.4]
  wire  storesToCheck_5_7; // @[LoadQueue.scala 131:10:@9649.4]
  wire  _T_8990; // @[LoadQueue.scala 131:81:@9652.4]
  wire  _T_8991; // @[LoadQueue.scala 131:72:@9653.4]
  wire  _T_8993; // @[LoadQueue.scala 132:33:@9654.4]
  wire  _T_8996; // @[LoadQueue.scala 132:41:@9656.4]
  wire  _T_8998; // @[LoadQueue.scala 132:9:@9657.4]
  wire  storesToCheck_5_8; // @[LoadQueue.scala 131:10:@9658.4]
  wire  _T_9004; // @[LoadQueue.scala 131:81:@9661.4]
  wire  _T_9005; // @[LoadQueue.scala 131:72:@9662.4]
  wire  _T_9007; // @[LoadQueue.scala 132:33:@9663.4]
  wire  _T_9010; // @[LoadQueue.scala 132:41:@9665.4]
  wire  _T_9012; // @[LoadQueue.scala 132:9:@9666.4]
  wire  storesToCheck_5_9; // @[LoadQueue.scala 131:10:@9667.4]
  wire  _T_9018; // @[LoadQueue.scala 131:81:@9670.4]
  wire  _T_9019; // @[LoadQueue.scala 131:72:@9671.4]
  wire  _T_9021; // @[LoadQueue.scala 132:33:@9672.4]
  wire  _T_9024; // @[LoadQueue.scala 132:41:@9674.4]
  wire  _T_9026; // @[LoadQueue.scala 132:9:@9675.4]
  wire  storesToCheck_5_10; // @[LoadQueue.scala 131:10:@9676.4]
  wire  _T_9032; // @[LoadQueue.scala 131:81:@9679.4]
  wire  _T_9033; // @[LoadQueue.scala 131:72:@9680.4]
  wire  _T_9035; // @[LoadQueue.scala 132:33:@9681.4]
  wire  _T_9038; // @[LoadQueue.scala 132:41:@9683.4]
  wire  _T_9040; // @[LoadQueue.scala 132:9:@9684.4]
  wire  storesToCheck_5_11; // @[LoadQueue.scala 131:10:@9685.4]
  wire  _T_9046; // @[LoadQueue.scala 131:81:@9688.4]
  wire  _T_9047; // @[LoadQueue.scala 131:72:@9689.4]
  wire  _T_9049; // @[LoadQueue.scala 132:33:@9690.4]
  wire  _T_9052; // @[LoadQueue.scala 132:41:@9692.4]
  wire  _T_9054; // @[LoadQueue.scala 132:9:@9693.4]
  wire  storesToCheck_5_12; // @[LoadQueue.scala 131:10:@9694.4]
  wire  _T_9060; // @[LoadQueue.scala 131:81:@9697.4]
  wire  _T_9061; // @[LoadQueue.scala 131:72:@9698.4]
  wire  _T_9063; // @[LoadQueue.scala 132:33:@9699.4]
  wire  _T_9066; // @[LoadQueue.scala 132:41:@9701.4]
  wire  _T_9068; // @[LoadQueue.scala 132:9:@9702.4]
  wire  storesToCheck_5_13; // @[LoadQueue.scala 131:10:@9703.4]
  wire  _T_9074; // @[LoadQueue.scala 131:81:@9706.4]
  wire  _T_9075; // @[LoadQueue.scala 131:72:@9707.4]
  wire  _T_9077; // @[LoadQueue.scala 132:33:@9708.4]
  wire  _T_9080; // @[LoadQueue.scala 132:41:@9710.4]
  wire  _T_9082; // @[LoadQueue.scala 132:9:@9711.4]
  wire  storesToCheck_5_14; // @[LoadQueue.scala 131:10:@9712.4]
  wire  _T_9088; // @[LoadQueue.scala 131:81:@9715.4]
  wire  storesToCheck_5_15; // @[LoadQueue.scala 131:10:@9721.4]
  wire  storesToCheck_6_0; // @[LoadQueue.scala 131:10:@9763.4]
  wire  _T_9138; // @[LoadQueue.scala 131:81:@9766.4]
  wire  _T_9139; // @[LoadQueue.scala 131:72:@9767.4]
  wire  _T_9141; // @[LoadQueue.scala 132:33:@9768.4]
  wire  _T_9144; // @[LoadQueue.scala 132:41:@9770.4]
  wire  _T_9146; // @[LoadQueue.scala 132:9:@9771.4]
  wire  storesToCheck_6_1; // @[LoadQueue.scala 131:10:@9772.4]
  wire  _T_9152; // @[LoadQueue.scala 131:81:@9775.4]
  wire  _T_9153; // @[LoadQueue.scala 131:72:@9776.4]
  wire  _T_9155; // @[LoadQueue.scala 132:33:@9777.4]
  wire  _T_9158; // @[LoadQueue.scala 132:41:@9779.4]
  wire  _T_9160; // @[LoadQueue.scala 132:9:@9780.4]
  wire  storesToCheck_6_2; // @[LoadQueue.scala 131:10:@9781.4]
  wire  _T_9166; // @[LoadQueue.scala 131:81:@9784.4]
  wire  _T_9167; // @[LoadQueue.scala 131:72:@9785.4]
  wire  _T_9169; // @[LoadQueue.scala 132:33:@9786.4]
  wire  _T_9172; // @[LoadQueue.scala 132:41:@9788.4]
  wire  _T_9174; // @[LoadQueue.scala 132:9:@9789.4]
  wire  storesToCheck_6_3; // @[LoadQueue.scala 131:10:@9790.4]
  wire  _T_9180; // @[LoadQueue.scala 131:81:@9793.4]
  wire  _T_9181; // @[LoadQueue.scala 131:72:@9794.4]
  wire  _T_9183; // @[LoadQueue.scala 132:33:@9795.4]
  wire  _T_9186; // @[LoadQueue.scala 132:41:@9797.4]
  wire  _T_9188; // @[LoadQueue.scala 132:9:@9798.4]
  wire  storesToCheck_6_4; // @[LoadQueue.scala 131:10:@9799.4]
  wire  _T_9194; // @[LoadQueue.scala 131:81:@9802.4]
  wire  _T_9195; // @[LoadQueue.scala 131:72:@9803.4]
  wire  _T_9197; // @[LoadQueue.scala 132:33:@9804.4]
  wire  _T_9200; // @[LoadQueue.scala 132:41:@9806.4]
  wire  _T_9202; // @[LoadQueue.scala 132:9:@9807.4]
  wire  storesToCheck_6_5; // @[LoadQueue.scala 131:10:@9808.4]
  wire  _T_9208; // @[LoadQueue.scala 131:81:@9811.4]
  wire  _T_9209; // @[LoadQueue.scala 131:72:@9812.4]
  wire  _T_9211; // @[LoadQueue.scala 132:33:@9813.4]
  wire  _T_9214; // @[LoadQueue.scala 132:41:@9815.4]
  wire  _T_9216; // @[LoadQueue.scala 132:9:@9816.4]
  wire  storesToCheck_6_6; // @[LoadQueue.scala 131:10:@9817.4]
  wire  _T_9222; // @[LoadQueue.scala 131:81:@9820.4]
  wire  _T_9223; // @[LoadQueue.scala 131:72:@9821.4]
  wire  _T_9225; // @[LoadQueue.scala 132:33:@9822.4]
  wire  _T_9228; // @[LoadQueue.scala 132:41:@9824.4]
  wire  _T_9230; // @[LoadQueue.scala 132:9:@9825.4]
  wire  storesToCheck_6_7; // @[LoadQueue.scala 131:10:@9826.4]
  wire  _T_9236; // @[LoadQueue.scala 131:81:@9829.4]
  wire  _T_9237; // @[LoadQueue.scala 131:72:@9830.4]
  wire  _T_9239; // @[LoadQueue.scala 132:33:@9831.4]
  wire  _T_9242; // @[LoadQueue.scala 132:41:@9833.4]
  wire  _T_9244; // @[LoadQueue.scala 132:9:@9834.4]
  wire  storesToCheck_6_8; // @[LoadQueue.scala 131:10:@9835.4]
  wire  _T_9250; // @[LoadQueue.scala 131:81:@9838.4]
  wire  _T_9251; // @[LoadQueue.scala 131:72:@9839.4]
  wire  _T_9253; // @[LoadQueue.scala 132:33:@9840.4]
  wire  _T_9256; // @[LoadQueue.scala 132:41:@9842.4]
  wire  _T_9258; // @[LoadQueue.scala 132:9:@9843.4]
  wire  storesToCheck_6_9; // @[LoadQueue.scala 131:10:@9844.4]
  wire  _T_9264; // @[LoadQueue.scala 131:81:@9847.4]
  wire  _T_9265; // @[LoadQueue.scala 131:72:@9848.4]
  wire  _T_9267; // @[LoadQueue.scala 132:33:@9849.4]
  wire  _T_9270; // @[LoadQueue.scala 132:41:@9851.4]
  wire  _T_9272; // @[LoadQueue.scala 132:9:@9852.4]
  wire  storesToCheck_6_10; // @[LoadQueue.scala 131:10:@9853.4]
  wire  _T_9278; // @[LoadQueue.scala 131:81:@9856.4]
  wire  _T_9279; // @[LoadQueue.scala 131:72:@9857.4]
  wire  _T_9281; // @[LoadQueue.scala 132:33:@9858.4]
  wire  _T_9284; // @[LoadQueue.scala 132:41:@9860.4]
  wire  _T_9286; // @[LoadQueue.scala 132:9:@9861.4]
  wire  storesToCheck_6_11; // @[LoadQueue.scala 131:10:@9862.4]
  wire  _T_9292; // @[LoadQueue.scala 131:81:@9865.4]
  wire  _T_9293; // @[LoadQueue.scala 131:72:@9866.4]
  wire  _T_9295; // @[LoadQueue.scala 132:33:@9867.4]
  wire  _T_9298; // @[LoadQueue.scala 132:41:@9869.4]
  wire  _T_9300; // @[LoadQueue.scala 132:9:@9870.4]
  wire  storesToCheck_6_12; // @[LoadQueue.scala 131:10:@9871.4]
  wire  _T_9306; // @[LoadQueue.scala 131:81:@9874.4]
  wire  _T_9307; // @[LoadQueue.scala 131:72:@9875.4]
  wire  _T_9309; // @[LoadQueue.scala 132:33:@9876.4]
  wire  _T_9312; // @[LoadQueue.scala 132:41:@9878.4]
  wire  _T_9314; // @[LoadQueue.scala 132:9:@9879.4]
  wire  storesToCheck_6_13; // @[LoadQueue.scala 131:10:@9880.4]
  wire  _T_9320; // @[LoadQueue.scala 131:81:@9883.4]
  wire  _T_9321; // @[LoadQueue.scala 131:72:@9884.4]
  wire  _T_9323; // @[LoadQueue.scala 132:33:@9885.4]
  wire  _T_9326; // @[LoadQueue.scala 132:41:@9887.4]
  wire  _T_9328; // @[LoadQueue.scala 132:9:@9888.4]
  wire  storesToCheck_6_14; // @[LoadQueue.scala 131:10:@9889.4]
  wire  _T_9334; // @[LoadQueue.scala 131:81:@9892.4]
  wire  storesToCheck_6_15; // @[LoadQueue.scala 131:10:@9898.4]
  wire  storesToCheck_7_0; // @[LoadQueue.scala 131:10:@9940.4]
  wire  _T_9384; // @[LoadQueue.scala 131:81:@9943.4]
  wire  _T_9385; // @[LoadQueue.scala 131:72:@9944.4]
  wire  _T_9387; // @[LoadQueue.scala 132:33:@9945.4]
  wire  _T_9390; // @[LoadQueue.scala 132:41:@9947.4]
  wire  _T_9392; // @[LoadQueue.scala 132:9:@9948.4]
  wire  storesToCheck_7_1; // @[LoadQueue.scala 131:10:@9949.4]
  wire  _T_9398; // @[LoadQueue.scala 131:81:@9952.4]
  wire  _T_9399; // @[LoadQueue.scala 131:72:@9953.4]
  wire  _T_9401; // @[LoadQueue.scala 132:33:@9954.4]
  wire  _T_9404; // @[LoadQueue.scala 132:41:@9956.4]
  wire  _T_9406; // @[LoadQueue.scala 132:9:@9957.4]
  wire  storesToCheck_7_2; // @[LoadQueue.scala 131:10:@9958.4]
  wire  _T_9412; // @[LoadQueue.scala 131:81:@9961.4]
  wire  _T_9413; // @[LoadQueue.scala 131:72:@9962.4]
  wire  _T_9415; // @[LoadQueue.scala 132:33:@9963.4]
  wire  _T_9418; // @[LoadQueue.scala 132:41:@9965.4]
  wire  _T_9420; // @[LoadQueue.scala 132:9:@9966.4]
  wire  storesToCheck_7_3; // @[LoadQueue.scala 131:10:@9967.4]
  wire  _T_9426; // @[LoadQueue.scala 131:81:@9970.4]
  wire  _T_9427; // @[LoadQueue.scala 131:72:@9971.4]
  wire  _T_9429; // @[LoadQueue.scala 132:33:@9972.4]
  wire  _T_9432; // @[LoadQueue.scala 132:41:@9974.4]
  wire  _T_9434; // @[LoadQueue.scala 132:9:@9975.4]
  wire  storesToCheck_7_4; // @[LoadQueue.scala 131:10:@9976.4]
  wire  _T_9440; // @[LoadQueue.scala 131:81:@9979.4]
  wire  _T_9441; // @[LoadQueue.scala 131:72:@9980.4]
  wire  _T_9443; // @[LoadQueue.scala 132:33:@9981.4]
  wire  _T_9446; // @[LoadQueue.scala 132:41:@9983.4]
  wire  _T_9448; // @[LoadQueue.scala 132:9:@9984.4]
  wire  storesToCheck_7_5; // @[LoadQueue.scala 131:10:@9985.4]
  wire  _T_9454; // @[LoadQueue.scala 131:81:@9988.4]
  wire  _T_9455; // @[LoadQueue.scala 131:72:@9989.4]
  wire  _T_9457; // @[LoadQueue.scala 132:33:@9990.4]
  wire  _T_9460; // @[LoadQueue.scala 132:41:@9992.4]
  wire  _T_9462; // @[LoadQueue.scala 132:9:@9993.4]
  wire  storesToCheck_7_6; // @[LoadQueue.scala 131:10:@9994.4]
  wire  _T_9468; // @[LoadQueue.scala 131:81:@9997.4]
  wire  _T_9469; // @[LoadQueue.scala 131:72:@9998.4]
  wire  _T_9471; // @[LoadQueue.scala 132:33:@9999.4]
  wire  _T_9474; // @[LoadQueue.scala 132:41:@10001.4]
  wire  _T_9476; // @[LoadQueue.scala 132:9:@10002.4]
  wire  storesToCheck_7_7; // @[LoadQueue.scala 131:10:@10003.4]
  wire  _T_9482; // @[LoadQueue.scala 131:81:@10006.4]
  wire  _T_9483; // @[LoadQueue.scala 131:72:@10007.4]
  wire  _T_9485; // @[LoadQueue.scala 132:33:@10008.4]
  wire  _T_9488; // @[LoadQueue.scala 132:41:@10010.4]
  wire  _T_9490; // @[LoadQueue.scala 132:9:@10011.4]
  wire  storesToCheck_7_8; // @[LoadQueue.scala 131:10:@10012.4]
  wire  _T_9496; // @[LoadQueue.scala 131:81:@10015.4]
  wire  _T_9497; // @[LoadQueue.scala 131:72:@10016.4]
  wire  _T_9499; // @[LoadQueue.scala 132:33:@10017.4]
  wire  _T_9502; // @[LoadQueue.scala 132:41:@10019.4]
  wire  _T_9504; // @[LoadQueue.scala 132:9:@10020.4]
  wire  storesToCheck_7_9; // @[LoadQueue.scala 131:10:@10021.4]
  wire  _T_9510; // @[LoadQueue.scala 131:81:@10024.4]
  wire  _T_9511; // @[LoadQueue.scala 131:72:@10025.4]
  wire  _T_9513; // @[LoadQueue.scala 132:33:@10026.4]
  wire  _T_9516; // @[LoadQueue.scala 132:41:@10028.4]
  wire  _T_9518; // @[LoadQueue.scala 132:9:@10029.4]
  wire  storesToCheck_7_10; // @[LoadQueue.scala 131:10:@10030.4]
  wire  _T_9524; // @[LoadQueue.scala 131:81:@10033.4]
  wire  _T_9525; // @[LoadQueue.scala 131:72:@10034.4]
  wire  _T_9527; // @[LoadQueue.scala 132:33:@10035.4]
  wire  _T_9530; // @[LoadQueue.scala 132:41:@10037.4]
  wire  _T_9532; // @[LoadQueue.scala 132:9:@10038.4]
  wire  storesToCheck_7_11; // @[LoadQueue.scala 131:10:@10039.4]
  wire  _T_9538; // @[LoadQueue.scala 131:81:@10042.4]
  wire  _T_9539; // @[LoadQueue.scala 131:72:@10043.4]
  wire  _T_9541; // @[LoadQueue.scala 132:33:@10044.4]
  wire  _T_9544; // @[LoadQueue.scala 132:41:@10046.4]
  wire  _T_9546; // @[LoadQueue.scala 132:9:@10047.4]
  wire  storesToCheck_7_12; // @[LoadQueue.scala 131:10:@10048.4]
  wire  _T_9552; // @[LoadQueue.scala 131:81:@10051.4]
  wire  _T_9553; // @[LoadQueue.scala 131:72:@10052.4]
  wire  _T_9555; // @[LoadQueue.scala 132:33:@10053.4]
  wire  _T_9558; // @[LoadQueue.scala 132:41:@10055.4]
  wire  _T_9560; // @[LoadQueue.scala 132:9:@10056.4]
  wire  storesToCheck_7_13; // @[LoadQueue.scala 131:10:@10057.4]
  wire  _T_9566; // @[LoadQueue.scala 131:81:@10060.4]
  wire  _T_9567; // @[LoadQueue.scala 131:72:@10061.4]
  wire  _T_9569; // @[LoadQueue.scala 132:33:@10062.4]
  wire  _T_9572; // @[LoadQueue.scala 132:41:@10064.4]
  wire  _T_9574; // @[LoadQueue.scala 132:9:@10065.4]
  wire  storesToCheck_7_14; // @[LoadQueue.scala 131:10:@10066.4]
  wire  _T_9580; // @[LoadQueue.scala 131:81:@10069.4]
  wire  storesToCheck_7_15; // @[LoadQueue.scala 131:10:@10075.4]
  wire  storesToCheck_8_0; // @[LoadQueue.scala 131:10:@10117.4]
  wire  _T_9630; // @[LoadQueue.scala 131:81:@10120.4]
  wire  _T_9631; // @[LoadQueue.scala 131:72:@10121.4]
  wire  _T_9633; // @[LoadQueue.scala 132:33:@10122.4]
  wire  _T_9636; // @[LoadQueue.scala 132:41:@10124.4]
  wire  _T_9638; // @[LoadQueue.scala 132:9:@10125.4]
  wire  storesToCheck_8_1; // @[LoadQueue.scala 131:10:@10126.4]
  wire  _T_9644; // @[LoadQueue.scala 131:81:@10129.4]
  wire  _T_9645; // @[LoadQueue.scala 131:72:@10130.4]
  wire  _T_9647; // @[LoadQueue.scala 132:33:@10131.4]
  wire  _T_9650; // @[LoadQueue.scala 132:41:@10133.4]
  wire  _T_9652; // @[LoadQueue.scala 132:9:@10134.4]
  wire  storesToCheck_8_2; // @[LoadQueue.scala 131:10:@10135.4]
  wire  _T_9658; // @[LoadQueue.scala 131:81:@10138.4]
  wire  _T_9659; // @[LoadQueue.scala 131:72:@10139.4]
  wire  _T_9661; // @[LoadQueue.scala 132:33:@10140.4]
  wire  _T_9664; // @[LoadQueue.scala 132:41:@10142.4]
  wire  _T_9666; // @[LoadQueue.scala 132:9:@10143.4]
  wire  storesToCheck_8_3; // @[LoadQueue.scala 131:10:@10144.4]
  wire  _T_9672; // @[LoadQueue.scala 131:81:@10147.4]
  wire  _T_9673; // @[LoadQueue.scala 131:72:@10148.4]
  wire  _T_9675; // @[LoadQueue.scala 132:33:@10149.4]
  wire  _T_9678; // @[LoadQueue.scala 132:41:@10151.4]
  wire  _T_9680; // @[LoadQueue.scala 132:9:@10152.4]
  wire  storesToCheck_8_4; // @[LoadQueue.scala 131:10:@10153.4]
  wire  _T_9686; // @[LoadQueue.scala 131:81:@10156.4]
  wire  _T_9687; // @[LoadQueue.scala 131:72:@10157.4]
  wire  _T_9689; // @[LoadQueue.scala 132:33:@10158.4]
  wire  _T_9692; // @[LoadQueue.scala 132:41:@10160.4]
  wire  _T_9694; // @[LoadQueue.scala 132:9:@10161.4]
  wire  storesToCheck_8_5; // @[LoadQueue.scala 131:10:@10162.4]
  wire  _T_9700; // @[LoadQueue.scala 131:81:@10165.4]
  wire  _T_9701; // @[LoadQueue.scala 131:72:@10166.4]
  wire  _T_9703; // @[LoadQueue.scala 132:33:@10167.4]
  wire  _T_9706; // @[LoadQueue.scala 132:41:@10169.4]
  wire  _T_9708; // @[LoadQueue.scala 132:9:@10170.4]
  wire  storesToCheck_8_6; // @[LoadQueue.scala 131:10:@10171.4]
  wire  _T_9714; // @[LoadQueue.scala 131:81:@10174.4]
  wire  _T_9715; // @[LoadQueue.scala 131:72:@10175.4]
  wire  _T_9717; // @[LoadQueue.scala 132:33:@10176.4]
  wire  _T_9720; // @[LoadQueue.scala 132:41:@10178.4]
  wire  _T_9722; // @[LoadQueue.scala 132:9:@10179.4]
  wire  storesToCheck_8_7; // @[LoadQueue.scala 131:10:@10180.4]
  wire  _T_9728; // @[LoadQueue.scala 131:81:@10183.4]
  wire  _T_9729; // @[LoadQueue.scala 131:72:@10184.4]
  wire  _T_9731; // @[LoadQueue.scala 132:33:@10185.4]
  wire  _T_9734; // @[LoadQueue.scala 132:41:@10187.4]
  wire  _T_9736; // @[LoadQueue.scala 132:9:@10188.4]
  wire  storesToCheck_8_8; // @[LoadQueue.scala 131:10:@10189.4]
  wire  _T_9742; // @[LoadQueue.scala 131:81:@10192.4]
  wire  _T_9743; // @[LoadQueue.scala 131:72:@10193.4]
  wire  _T_9745; // @[LoadQueue.scala 132:33:@10194.4]
  wire  _T_9748; // @[LoadQueue.scala 132:41:@10196.4]
  wire  _T_9750; // @[LoadQueue.scala 132:9:@10197.4]
  wire  storesToCheck_8_9; // @[LoadQueue.scala 131:10:@10198.4]
  wire  _T_9756; // @[LoadQueue.scala 131:81:@10201.4]
  wire  _T_9757; // @[LoadQueue.scala 131:72:@10202.4]
  wire  _T_9759; // @[LoadQueue.scala 132:33:@10203.4]
  wire  _T_9762; // @[LoadQueue.scala 132:41:@10205.4]
  wire  _T_9764; // @[LoadQueue.scala 132:9:@10206.4]
  wire  storesToCheck_8_10; // @[LoadQueue.scala 131:10:@10207.4]
  wire  _T_9770; // @[LoadQueue.scala 131:81:@10210.4]
  wire  _T_9771; // @[LoadQueue.scala 131:72:@10211.4]
  wire  _T_9773; // @[LoadQueue.scala 132:33:@10212.4]
  wire  _T_9776; // @[LoadQueue.scala 132:41:@10214.4]
  wire  _T_9778; // @[LoadQueue.scala 132:9:@10215.4]
  wire  storesToCheck_8_11; // @[LoadQueue.scala 131:10:@10216.4]
  wire  _T_9784; // @[LoadQueue.scala 131:81:@10219.4]
  wire  _T_9785; // @[LoadQueue.scala 131:72:@10220.4]
  wire  _T_9787; // @[LoadQueue.scala 132:33:@10221.4]
  wire  _T_9790; // @[LoadQueue.scala 132:41:@10223.4]
  wire  _T_9792; // @[LoadQueue.scala 132:9:@10224.4]
  wire  storesToCheck_8_12; // @[LoadQueue.scala 131:10:@10225.4]
  wire  _T_9798; // @[LoadQueue.scala 131:81:@10228.4]
  wire  _T_9799; // @[LoadQueue.scala 131:72:@10229.4]
  wire  _T_9801; // @[LoadQueue.scala 132:33:@10230.4]
  wire  _T_9804; // @[LoadQueue.scala 132:41:@10232.4]
  wire  _T_9806; // @[LoadQueue.scala 132:9:@10233.4]
  wire  storesToCheck_8_13; // @[LoadQueue.scala 131:10:@10234.4]
  wire  _T_9812; // @[LoadQueue.scala 131:81:@10237.4]
  wire  _T_9813; // @[LoadQueue.scala 131:72:@10238.4]
  wire  _T_9815; // @[LoadQueue.scala 132:33:@10239.4]
  wire  _T_9818; // @[LoadQueue.scala 132:41:@10241.4]
  wire  _T_9820; // @[LoadQueue.scala 132:9:@10242.4]
  wire  storesToCheck_8_14; // @[LoadQueue.scala 131:10:@10243.4]
  wire  _T_9826; // @[LoadQueue.scala 131:81:@10246.4]
  wire  storesToCheck_8_15; // @[LoadQueue.scala 131:10:@10252.4]
  wire  storesToCheck_9_0; // @[LoadQueue.scala 131:10:@10294.4]
  wire  _T_9876; // @[LoadQueue.scala 131:81:@10297.4]
  wire  _T_9877; // @[LoadQueue.scala 131:72:@10298.4]
  wire  _T_9879; // @[LoadQueue.scala 132:33:@10299.4]
  wire  _T_9882; // @[LoadQueue.scala 132:41:@10301.4]
  wire  _T_9884; // @[LoadQueue.scala 132:9:@10302.4]
  wire  storesToCheck_9_1; // @[LoadQueue.scala 131:10:@10303.4]
  wire  _T_9890; // @[LoadQueue.scala 131:81:@10306.4]
  wire  _T_9891; // @[LoadQueue.scala 131:72:@10307.4]
  wire  _T_9893; // @[LoadQueue.scala 132:33:@10308.4]
  wire  _T_9896; // @[LoadQueue.scala 132:41:@10310.4]
  wire  _T_9898; // @[LoadQueue.scala 132:9:@10311.4]
  wire  storesToCheck_9_2; // @[LoadQueue.scala 131:10:@10312.4]
  wire  _T_9904; // @[LoadQueue.scala 131:81:@10315.4]
  wire  _T_9905; // @[LoadQueue.scala 131:72:@10316.4]
  wire  _T_9907; // @[LoadQueue.scala 132:33:@10317.4]
  wire  _T_9910; // @[LoadQueue.scala 132:41:@10319.4]
  wire  _T_9912; // @[LoadQueue.scala 132:9:@10320.4]
  wire  storesToCheck_9_3; // @[LoadQueue.scala 131:10:@10321.4]
  wire  _T_9918; // @[LoadQueue.scala 131:81:@10324.4]
  wire  _T_9919; // @[LoadQueue.scala 131:72:@10325.4]
  wire  _T_9921; // @[LoadQueue.scala 132:33:@10326.4]
  wire  _T_9924; // @[LoadQueue.scala 132:41:@10328.4]
  wire  _T_9926; // @[LoadQueue.scala 132:9:@10329.4]
  wire  storesToCheck_9_4; // @[LoadQueue.scala 131:10:@10330.4]
  wire  _T_9932; // @[LoadQueue.scala 131:81:@10333.4]
  wire  _T_9933; // @[LoadQueue.scala 131:72:@10334.4]
  wire  _T_9935; // @[LoadQueue.scala 132:33:@10335.4]
  wire  _T_9938; // @[LoadQueue.scala 132:41:@10337.4]
  wire  _T_9940; // @[LoadQueue.scala 132:9:@10338.4]
  wire  storesToCheck_9_5; // @[LoadQueue.scala 131:10:@10339.4]
  wire  _T_9946; // @[LoadQueue.scala 131:81:@10342.4]
  wire  _T_9947; // @[LoadQueue.scala 131:72:@10343.4]
  wire  _T_9949; // @[LoadQueue.scala 132:33:@10344.4]
  wire  _T_9952; // @[LoadQueue.scala 132:41:@10346.4]
  wire  _T_9954; // @[LoadQueue.scala 132:9:@10347.4]
  wire  storesToCheck_9_6; // @[LoadQueue.scala 131:10:@10348.4]
  wire  _T_9960; // @[LoadQueue.scala 131:81:@10351.4]
  wire  _T_9961; // @[LoadQueue.scala 131:72:@10352.4]
  wire  _T_9963; // @[LoadQueue.scala 132:33:@10353.4]
  wire  _T_9966; // @[LoadQueue.scala 132:41:@10355.4]
  wire  _T_9968; // @[LoadQueue.scala 132:9:@10356.4]
  wire  storesToCheck_9_7; // @[LoadQueue.scala 131:10:@10357.4]
  wire  _T_9974; // @[LoadQueue.scala 131:81:@10360.4]
  wire  _T_9975; // @[LoadQueue.scala 131:72:@10361.4]
  wire  _T_9977; // @[LoadQueue.scala 132:33:@10362.4]
  wire  _T_9980; // @[LoadQueue.scala 132:41:@10364.4]
  wire  _T_9982; // @[LoadQueue.scala 132:9:@10365.4]
  wire  storesToCheck_9_8; // @[LoadQueue.scala 131:10:@10366.4]
  wire  _T_9988; // @[LoadQueue.scala 131:81:@10369.4]
  wire  _T_9989; // @[LoadQueue.scala 131:72:@10370.4]
  wire  _T_9991; // @[LoadQueue.scala 132:33:@10371.4]
  wire  _T_9994; // @[LoadQueue.scala 132:41:@10373.4]
  wire  _T_9996; // @[LoadQueue.scala 132:9:@10374.4]
  wire  storesToCheck_9_9; // @[LoadQueue.scala 131:10:@10375.4]
  wire  _T_10002; // @[LoadQueue.scala 131:81:@10378.4]
  wire  _T_10003; // @[LoadQueue.scala 131:72:@10379.4]
  wire  _T_10005; // @[LoadQueue.scala 132:33:@10380.4]
  wire  _T_10008; // @[LoadQueue.scala 132:41:@10382.4]
  wire  _T_10010; // @[LoadQueue.scala 132:9:@10383.4]
  wire  storesToCheck_9_10; // @[LoadQueue.scala 131:10:@10384.4]
  wire  _T_10016; // @[LoadQueue.scala 131:81:@10387.4]
  wire  _T_10017; // @[LoadQueue.scala 131:72:@10388.4]
  wire  _T_10019; // @[LoadQueue.scala 132:33:@10389.4]
  wire  _T_10022; // @[LoadQueue.scala 132:41:@10391.4]
  wire  _T_10024; // @[LoadQueue.scala 132:9:@10392.4]
  wire  storesToCheck_9_11; // @[LoadQueue.scala 131:10:@10393.4]
  wire  _T_10030; // @[LoadQueue.scala 131:81:@10396.4]
  wire  _T_10031; // @[LoadQueue.scala 131:72:@10397.4]
  wire  _T_10033; // @[LoadQueue.scala 132:33:@10398.4]
  wire  _T_10036; // @[LoadQueue.scala 132:41:@10400.4]
  wire  _T_10038; // @[LoadQueue.scala 132:9:@10401.4]
  wire  storesToCheck_9_12; // @[LoadQueue.scala 131:10:@10402.4]
  wire  _T_10044; // @[LoadQueue.scala 131:81:@10405.4]
  wire  _T_10045; // @[LoadQueue.scala 131:72:@10406.4]
  wire  _T_10047; // @[LoadQueue.scala 132:33:@10407.4]
  wire  _T_10050; // @[LoadQueue.scala 132:41:@10409.4]
  wire  _T_10052; // @[LoadQueue.scala 132:9:@10410.4]
  wire  storesToCheck_9_13; // @[LoadQueue.scala 131:10:@10411.4]
  wire  _T_10058; // @[LoadQueue.scala 131:81:@10414.4]
  wire  _T_10059; // @[LoadQueue.scala 131:72:@10415.4]
  wire  _T_10061; // @[LoadQueue.scala 132:33:@10416.4]
  wire  _T_10064; // @[LoadQueue.scala 132:41:@10418.4]
  wire  _T_10066; // @[LoadQueue.scala 132:9:@10419.4]
  wire  storesToCheck_9_14; // @[LoadQueue.scala 131:10:@10420.4]
  wire  _T_10072; // @[LoadQueue.scala 131:81:@10423.4]
  wire  storesToCheck_9_15; // @[LoadQueue.scala 131:10:@10429.4]
  wire  storesToCheck_10_0; // @[LoadQueue.scala 131:10:@10471.4]
  wire  _T_10122; // @[LoadQueue.scala 131:81:@10474.4]
  wire  _T_10123; // @[LoadQueue.scala 131:72:@10475.4]
  wire  _T_10125; // @[LoadQueue.scala 132:33:@10476.4]
  wire  _T_10128; // @[LoadQueue.scala 132:41:@10478.4]
  wire  _T_10130; // @[LoadQueue.scala 132:9:@10479.4]
  wire  storesToCheck_10_1; // @[LoadQueue.scala 131:10:@10480.4]
  wire  _T_10136; // @[LoadQueue.scala 131:81:@10483.4]
  wire  _T_10137; // @[LoadQueue.scala 131:72:@10484.4]
  wire  _T_10139; // @[LoadQueue.scala 132:33:@10485.4]
  wire  _T_10142; // @[LoadQueue.scala 132:41:@10487.4]
  wire  _T_10144; // @[LoadQueue.scala 132:9:@10488.4]
  wire  storesToCheck_10_2; // @[LoadQueue.scala 131:10:@10489.4]
  wire  _T_10150; // @[LoadQueue.scala 131:81:@10492.4]
  wire  _T_10151; // @[LoadQueue.scala 131:72:@10493.4]
  wire  _T_10153; // @[LoadQueue.scala 132:33:@10494.4]
  wire  _T_10156; // @[LoadQueue.scala 132:41:@10496.4]
  wire  _T_10158; // @[LoadQueue.scala 132:9:@10497.4]
  wire  storesToCheck_10_3; // @[LoadQueue.scala 131:10:@10498.4]
  wire  _T_10164; // @[LoadQueue.scala 131:81:@10501.4]
  wire  _T_10165; // @[LoadQueue.scala 131:72:@10502.4]
  wire  _T_10167; // @[LoadQueue.scala 132:33:@10503.4]
  wire  _T_10170; // @[LoadQueue.scala 132:41:@10505.4]
  wire  _T_10172; // @[LoadQueue.scala 132:9:@10506.4]
  wire  storesToCheck_10_4; // @[LoadQueue.scala 131:10:@10507.4]
  wire  _T_10178; // @[LoadQueue.scala 131:81:@10510.4]
  wire  _T_10179; // @[LoadQueue.scala 131:72:@10511.4]
  wire  _T_10181; // @[LoadQueue.scala 132:33:@10512.4]
  wire  _T_10184; // @[LoadQueue.scala 132:41:@10514.4]
  wire  _T_10186; // @[LoadQueue.scala 132:9:@10515.4]
  wire  storesToCheck_10_5; // @[LoadQueue.scala 131:10:@10516.4]
  wire  _T_10192; // @[LoadQueue.scala 131:81:@10519.4]
  wire  _T_10193; // @[LoadQueue.scala 131:72:@10520.4]
  wire  _T_10195; // @[LoadQueue.scala 132:33:@10521.4]
  wire  _T_10198; // @[LoadQueue.scala 132:41:@10523.4]
  wire  _T_10200; // @[LoadQueue.scala 132:9:@10524.4]
  wire  storesToCheck_10_6; // @[LoadQueue.scala 131:10:@10525.4]
  wire  _T_10206; // @[LoadQueue.scala 131:81:@10528.4]
  wire  _T_10207; // @[LoadQueue.scala 131:72:@10529.4]
  wire  _T_10209; // @[LoadQueue.scala 132:33:@10530.4]
  wire  _T_10212; // @[LoadQueue.scala 132:41:@10532.4]
  wire  _T_10214; // @[LoadQueue.scala 132:9:@10533.4]
  wire  storesToCheck_10_7; // @[LoadQueue.scala 131:10:@10534.4]
  wire  _T_10220; // @[LoadQueue.scala 131:81:@10537.4]
  wire  _T_10221; // @[LoadQueue.scala 131:72:@10538.4]
  wire  _T_10223; // @[LoadQueue.scala 132:33:@10539.4]
  wire  _T_10226; // @[LoadQueue.scala 132:41:@10541.4]
  wire  _T_10228; // @[LoadQueue.scala 132:9:@10542.4]
  wire  storesToCheck_10_8; // @[LoadQueue.scala 131:10:@10543.4]
  wire  _T_10234; // @[LoadQueue.scala 131:81:@10546.4]
  wire  _T_10235; // @[LoadQueue.scala 131:72:@10547.4]
  wire  _T_10237; // @[LoadQueue.scala 132:33:@10548.4]
  wire  _T_10240; // @[LoadQueue.scala 132:41:@10550.4]
  wire  _T_10242; // @[LoadQueue.scala 132:9:@10551.4]
  wire  storesToCheck_10_9; // @[LoadQueue.scala 131:10:@10552.4]
  wire  _T_10248; // @[LoadQueue.scala 131:81:@10555.4]
  wire  _T_10249; // @[LoadQueue.scala 131:72:@10556.4]
  wire  _T_10251; // @[LoadQueue.scala 132:33:@10557.4]
  wire  _T_10254; // @[LoadQueue.scala 132:41:@10559.4]
  wire  _T_10256; // @[LoadQueue.scala 132:9:@10560.4]
  wire  storesToCheck_10_10; // @[LoadQueue.scala 131:10:@10561.4]
  wire  _T_10262; // @[LoadQueue.scala 131:81:@10564.4]
  wire  _T_10263; // @[LoadQueue.scala 131:72:@10565.4]
  wire  _T_10265; // @[LoadQueue.scala 132:33:@10566.4]
  wire  _T_10268; // @[LoadQueue.scala 132:41:@10568.4]
  wire  _T_10270; // @[LoadQueue.scala 132:9:@10569.4]
  wire  storesToCheck_10_11; // @[LoadQueue.scala 131:10:@10570.4]
  wire  _T_10276; // @[LoadQueue.scala 131:81:@10573.4]
  wire  _T_10277; // @[LoadQueue.scala 131:72:@10574.4]
  wire  _T_10279; // @[LoadQueue.scala 132:33:@10575.4]
  wire  _T_10282; // @[LoadQueue.scala 132:41:@10577.4]
  wire  _T_10284; // @[LoadQueue.scala 132:9:@10578.4]
  wire  storesToCheck_10_12; // @[LoadQueue.scala 131:10:@10579.4]
  wire  _T_10290; // @[LoadQueue.scala 131:81:@10582.4]
  wire  _T_10291; // @[LoadQueue.scala 131:72:@10583.4]
  wire  _T_10293; // @[LoadQueue.scala 132:33:@10584.4]
  wire  _T_10296; // @[LoadQueue.scala 132:41:@10586.4]
  wire  _T_10298; // @[LoadQueue.scala 132:9:@10587.4]
  wire  storesToCheck_10_13; // @[LoadQueue.scala 131:10:@10588.4]
  wire  _T_10304; // @[LoadQueue.scala 131:81:@10591.4]
  wire  _T_10305; // @[LoadQueue.scala 131:72:@10592.4]
  wire  _T_10307; // @[LoadQueue.scala 132:33:@10593.4]
  wire  _T_10310; // @[LoadQueue.scala 132:41:@10595.4]
  wire  _T_10312; // @[LoadQueue.scala 132:9:@10596.4]
  wire  storesToCheck_10_14; // @[LoadQueue.scala 131:10:@10597.4]
  wire  _T_10318; // @[LoadQueue.scala 131:81:@10600.4]
  wire  storesToCheck_10_15; // @[LoadQueue.scala 131:10:@10606.4]
  wire  storesToCheck_11_0; // @[LoadQueue.scala 131:10:@10648.4]
  wire  _T_10368; // @[LoadQueue.scala 131:81:@10651.4]
  wire  _T_10369; // @[LoadQueue.scala 131:72:@10652.4]
  wire  _T_10371; // @[LoadQueue.scala 132:33:@10653.4]
  wire  _T_10374; // @[LoadQueue.scala 132:41:@10655.4]
  wire  _T_10376; // @[LoadQueue.scala 132:9:@10656.4]
  wire  storesToCheck_11_1; // @[LoadQueue.scala 131:10:@10657.4]
  wire  _T_10382; // @[LoadQueue.scala 131:81:@10660.4]
  wire  _T_10383; // @[LoadQueue.scala 131:72:@10661.4]
  wire  _T_10385; // @[LoadQueue.scala 132:33:@10662.4]
  wire  _T_10388; // @[LoadQueue.scala 132:41:@10664.4]
  wire  _T_10390; // @[LoadQueue.scala 132:9:@10665.4]
  wire  storesToCheck_11_2; // @[LoadQueue.scala 131:10:@10666.4]
  wire  _T_10396; // @[LoadQueue.scala 131:81:@10669.4]
  wire  _T_10397; // @[LoadQueue.scala 131:72:@10670.4]
  wire  _T_10399; // @[LoadQueue.scala 132:33:@10671.4]
  wire  _T_10402; // @[LoadQueue.scala 132:41:@10673.4]
  wire  _T_10404; // @[LoadQueue.scala 132:9:@10674.4]
  wire  storesToCheck_11_3; // @[LoadQueue.scala 131:10:@10675.4]
  wire  _T_10410; // @[LoadQueue.scala 131:81:@10678.4]
  wire  _T_10411; // @[LoadQueue.scala 131:72:@10679.4]
  wire  _T_10413; // @[LoadQueue.scala 132:33:@10680.4]
  wire  _T_10416; // @[LoadQueue.scala 132:41:@10682.4]
  wire  _T_10418; // @[LoadQueue.scala 132:9:@10683.4]
  wire  storesToCheck_11_4; // @[LoadQueue.scala 131:10:@10684.4]
  wire  _T_10424; // @[LoadQueue.scala 131:81:@10687.4]
  wire  _T_10425; // @[LoadQueue.scala 131:72:@10688.4]
  wire  _T_10427; // @[LoadQueue.scala 132:33:@10689.4]
  wire  _T_10430; // @[LoadQueue.scala 132:41:@10691.4]
  wire  _T_10432; // @[LoadQueue.scala 132:9:@10692.4]
  wire  storesToCheck_11_5; // @[LoadQueue.scala 131:10:@10693.4]
  wire  _T_10438; // @[LoadQueue.scala 131:81:@10696.4]
  wire  _T_10439; // @[LoadQueue.scala 131:72:@10697.4]
  wire  _T_10441; // @[LoadQueue.scala 132:33:@10698.4]
  wire  _T_10444; // @[LoadQueue.scala 132:41:@10700.4]
  wire  _T_10446; // @[LoadQueue.scala 132:9:@10701.4]
  wire  storesToCheck_11_6; // @[LoadQueue.scala 131:10:@10702.4]
  wire  _T_10452; // @[LoadQueue.scala 131:81:@10705.4]
  wire  _T_10453; // @[LoadQueue.scala 131:72:@10706.4]
  wire  _T_10455; // @[LoadQueue.scala 132:33:@10707.4]
  wire  _T_10458; // @[LoadQueue.scala 132:41:@10709.4]
  wire  _T_10460; // @[LoadQueue.scala 132:9:@10710.4]
  wire  storesToCheck_11_7; // @[LoadQueue.scala 131:10:@10711.4]
  wire  _T_10466; // @[LoadQueue.scala 131:81:@10714.4]
  wire  _T_10467; // @[LoadQueue.scala 131:72:@10715.4]
  wire  _T_10469; // @[LoadQueue.scala 132:33:@10716.4]
  wire  _T_10472; // @[LoadQueue.scala 132:41:@10718.4]
  wire  _T_10474; // @[LoadQueue.scala 132:9:@10719.4]
  wire  storesToCheck_11_8; // @[LoadQueue.scala 131:10:@10720.4]
  wire  _T_10480; // @[LoadQueue.scala 131:81:@10723.4]
  wire  _T_10481; // @[LoadQueue.scala 131:72:@10724.4]
  wire  _T_10483; // @[LoadQueue.scala 132:33:@10725.4]
  wire  _T_10486; // @[LoadQueue.scala 132:41:@10727.4]
  wire  _T_10488; // @[LoadQueue.scala 132:9:@10728.4]
  wire  storesToCheck_11_9; // @[LoadQueue.scala 131:10:@10729.4]
  wire  _T_10494; // @[LoadQueue.scala 131:81:@10732.4]
  wire  _T_10495; // @[LoadQueue.scala 131:72:@10733.4]
  wire  _T_10497; // @[LoadQueue.scala 132:33:@10734.4]
  wire  _T_10500; // @[LoadQueue.scala 132:41:@10736.4]
  wire  _T_10502; // @[LoadQueue.scala 132:9:@10737.4]
  wire  storesToCheck_11_10; // @[LoadQueue.scala 131:10:@10738.4]
  wire  _T_10508; // @[LoadQueue.scala 131:81:@10741.4]
  wire  _T_10509; // @[LoadQueue.scala 131:72:@10742.4]
  wire  _T_10511; // @[LoadQueue.scala 132:33:@10743.4]
  wire  _T_10514; // @[LoadQueue.scala 132:41:@10745.4]
  wire  _T_10516; // @[LoadQueue.scala 132:9:@10746.4]
  wire  storesToCheck_11_11; // @[LoadQueue.scala 131:10:@10747.4]
  wire  _T_10522; // @[LoadQueue.scala 131:81:@10750.4]
  wire  _T_10523; // @[LoadQueue.scala 131:72:@10751.4]
  wire  _T_10525; // @[LoadQueue.scala 132:33:@10752.4]
  wire  _T_10528; // @[LoadQueue.scala 132:41:@10754.4]
  wire  _T_10530; // @[LoadQueue.scala 132:9:@10755.4]
  wire  storesToCheck_11_12; // @[LoadQueue.scala 131:10:@10756.4]
  wire  _T_10536; // @[LoadQueue.scala 131:81:@10759.4]
  wire  _T_10537; // @[LoadQueue.scala 131:72:@10760.4]
  wire  _T_10539; // @[LoadQueue.scala 132:33:@10761.4]
  wire  _T_10542; // @[LoadQueue.scala 132:41:@10763.4]
  wire  _T_10544; // @[LoadQueue.scala 132:9:@10764.4]
  wire  storesToCheck_11_13; // @[LoadQueue.scala 131:10:@10765.4]
  wire  _T_10550; // @[LoadQueue.scala 131:81:@10768.4]
  wire  _T_10551; // @[LoadQueue.scala 131:72:@10769.4]
  wire  _T_10553; // @[LoadQueue.scala 132:33:@10770.4]
  wire  _T_10556; // @[LoadQueue.scala 132:41:@10772.4]
  wire  _T_10558; // @[LoadQueue.scala 132:9:@10773.4]
  wire  storesToCheck_11_14; // @[LoadQueue.scala 131:10:@10774.4]
  wire  _T_10564; // @[LoadQueue.scala 131:81:@10777.4]
  wire  storesToCheck_11_15; // @[LoadQueue.scala 131:10:@10783.4]
  wire  storesToCheck_12_0; // @[LoadQueue.scala 131:10:@10825.4]
  wire  _T_10614; // @[LoadQueue.scala 131:81:@10828.4]
  wire  _T_10615; // @[LoadQueue.scala 131:72:@10829.4]
  wire  _T_10617; // @[LoadQueue.scala 132:33:@10830.4]
  wire  _T_10620; // @[LoadQueue.scala 132:41:@10832.4]
  wire  _T_10622; // @[LoadQueue.scala 132:9:@10833.4]
  wire  storesToCheck_12_1; // @[LoadQueue.scala 131:10:@10834.4]
  wire  _T_10628; // @[LoadQueue.scala 131:81:@10837.4]
  wire  _T_10629; // @[LoadQueue.scala 131:72:@10838.4]
  wire  _T_10631; // @[LoadQueue.scala 132:33:@10839.4]
  wire  _T_10634; // @[LoadQueue.scala 132:41:@10841.4]
  wire  _T_10636; // @[LoadQueue.scala 132:9:@10842.4]
  wire  storesToCheck_12_2; // @[LoadQueue.scala 131:10:@10843.4]
  wire  _T_10642; // @[LoadQueue.scala 131:81:@10846.4]
  wire  _T_10643; // @[LoadQueue.scala 131:72:@10847.4]
  wire  _T_10645; // @[LoadQueue.scala 132:33:@10848.4]
  wire  _T_10648; // @[LoadQueue.scala 132:41:@10850.4]
  wire  _T_10650; // @[LoadQueue.scala 132:9:@10851.4]
  wire  storesToCheck_12_3; // @[LoadQueue.scala 131:10:@10852.4]
  wire  _T_10656; // @[LoadQueue.scala 131:81:@10855.4]
  wire  _T_10657; // @[LoadQueue.scala 131:72:@10856.4]
  wire  _T_10659; // @[LoadQueue.scala 132:33:@10857.4]
  wire  _T_10662; // @[LoadQueue.scala 132:41:@10859.4]
  wire  _T_10664; // @[LoadQueue.scala 132:9:@10860.4]
  wire  storesToCheck_12_4; // @[LoadQueue.scala 131:10:@10861.4]
  wire  _T_10670; // @[LoadQueue.scala 131:81:@10864.4]
  wire  _T_10671; // @[LoadQueue.scala 131:72:@10865.4]
  wire  _T_10673; // @[LoadQueue.scala 132:33:@10866.4]
  wire  _T_10676; // @[LoadQueue.scala 132:41:@10868.4]
  wire  _T_10678; // @[LoadQueue.scala 132:9:@10869.4]
  wire  storesToCheck_12_5; // @[LoadQueue.scala 131:10:@10870.4]
  wire  _T_10684; // @[LoadQueue.scala 131:81:@10873.4]
  wire  _T_10685; // @[LoadQueue.scala 131:72:@10874.4]
  wire  _T_10687; // @[LoadQueue.scala 132:33:@10875.4]
  wire  _T_10690; // @[LoadQueue.scala 132:41:@10877.4]
  wire  _T_10692; // @[LoadQueue.scala 132:9:@10878.4]
  wire  storesToCheck_12_6; // @[LoadQueue.scala 131:10:@10879.4]
  wire  _T_10698; // @[LoadQueue.scala 131:81:@10882.4]
  wire  _T_10699; // @[LoadQueue.scala 131:72:@10883.4]
  wire  _T_10701; // @[LoadQueue.scala 132:33:@10884.4]
  wire  _T_10704; // @[LoadQueue.scala 132:41:@10886.4]
  wire  _T_10706; // @[LoadQueue.scala 132:9:@10887.4]
  wire  storesToCheck_12_7; // @[LoadQueue.scala 131:10:@10888.4]
  wire  _T_10712; // @[LoadQueue.scala 131:81:@10891.4]
  wire  _T_10713; // @[LoadQueue.scala 131:72:@10892.4]
  wire  _T_10715; // @[LoadQueue.scala 132:33:@10893.4]
  wire  _T_10718; // @[LoadQueue.scala 132:41:@10895.4]
  wire  _T_10720; // @[LoadQueue.scala 132:9:@10896.4]
  wire  storesToCheck_12_8; // @[LoadQueue.scala 131:10:@10897.4]
  wire  _T_10726; // @[LoadQueue.scala 131:81:@10900.4]
  wire  _T_10727; // @[LoadQueue.scala 131:72:@10901.4]
  wire  _T_10729; // @[LoadQueue.scala 132:33:@10902.4]
  wire  _T_10732; // @[LoadQueue.scala 132:41:@10904.4]
  wire  _T_10734; // @[LoadQueue.scala 132:9:@10905.4]
  wire  storesToCheck_12_9; // @[LoadQueue.scala 131:10:@10906.4]
  wire  _T_10740; // @[LoadQueue.scala 131:81:@10909.4]
  wire  _T_10741; // @[LoadQueue.scala 131:72:@10910.4]
  wire  _T_10743; // @[LoadQueue.scala 132:33:@10911.4]
  wire  _T_10746; // @[LoadQueue.scala 132:41:@10913.4]
  wire  _T_10748; // @[LoadQueue.scala 132:9:@10914.4]
  wire  storesToCheck_12_10; // @[LoadQueue.scala 131:10:@10915.4]
  wire  _T_10754; // @[LoadQueue.scala 131:81:@10918.4]
  wire  _T_10755; // @[LoadQueue.scala 131:72:@10919.4]
  wire  _T_10757; // @[LoadQueue.scala 132:33:@10920.4]
  wire  _T_10760; // @[LoadQueue.scala 132:41:@10922.4]
  wire  _T_10762; // @[LoadQueue.scala 132:9:@10923.4]
  wire  storesToCheck_12_11; // @[LoadQueue.scala 131:10:@10924.4]
  wire  _T_10768; // @[LoadQueue.scala 131:81:@10927.4]
  wire  _T_10769; // @[LoadQueue.scala 131:72:@10928.4]
  wire  _T_10771; // @[LoadQueue.scala 132:33:@10929.4]
  wire  _T_10774; // @[LoadQueue.scala 132:41:@10931.4]
  wire  _T_10776; // @[LoadQueue.scala 132:9:@10932.4]
  wire  storesToCheck_12_12; // @[LoadQueue.scala 131:10:@10933.4]
  wire  _T_10782; // @[LoadQueue.scala 131:81:@10936.4]
  wire  _T_10783; // @[LoadQueue.scala 131:72:@10937.4]
  wire  _T_10785; // @[LoadQueue.scala 132:33:@10938.4]
  wire  _T_10788; // @[LoadQueue.scala 132:41:@10940.4]
  wire  _T_10790; // @[LoadQueue.scala 132:9:@10941.4]
  wire  storesToCheck_12_13; // @[LoadQueue.scala 131:10:@10942.4]
  wire  _T_10796; // @[LoadQueue.scala 131:81:@10945.4]
  wire  _T_10797; // @[LoadQueue.scala 131:72:@10946.4]
  wire  _T_10799; // @[LoadQueue.scala 132:33:@10947.4]
  wire  _T_10802; // @[LoadQueue.scala 132:41:@10949.4]
  wire  _T_10804; // @[LoadQueue.scala 132:9:@10950.4]
  wire  storesToCheck_12_14; // @[LoadQueue.scala 131:10:@10951.4]
  wire  _T_10810; // @[LoadQueue.scala 131:81:@10954.4]
  wire  storesToCheck_12_15; // @[LoadQueue.scala 131:10:@10960.4]
  wire  storesToCheck_13_0; // @[LoadQueue.scala 131:10:@11002.4]
  wire  _T_10860; // @[LoadQueue.scala 131:81:@11005.4]
  wire  _T_10861; // @[LoadQueue.scala 131:72:@11006.4]
  wire  _T_10863; // @[LoadQueue.scala 132:33:@11007.4]
  wire  _T_10866; // @[LoadQueue.scala 132:41:@11009.4]
  wire  _T_10868; // @[LoadQueue.scala 132:9:@11010.4]
  wire  storesToCheck_13_1; // @[LoadQueue.scala 131:10:@11011.4]
  wire  _T_10874; // @[LoadQueue.scala 131:81:@11014.4]
  wire  _T_10875; // @[LoadQueue.scala 131:72:@11015.4]
  wire  _T_10877; // @[LoadQueue.scala 132:33:@11016.4]
  wire  _T_10880; // @[LoadQueue.scala 132:41:@11018.4]
  wire  _T_10882; // @[LoadQueue.scala 132:9:@11019.4]
  wire  storesToCheck_13_2; // @[LoadQueue.scala 131:10:@11020.4]
  wire  _T_10888; // @[LoadQueue.scala 131:81:@11023.4]
  wire  _T_10889; // @[LoadQueue.scala 131:72:@11024.4]
  wire  _T_10891; // @[LoadQueue.scala 132:33:@11025.4]
  wire  _T_10894; // @[LoadQueue.scala 132:41:@11027.4]
  wire  _T_10896; // @[LoadQueue.scala 132:9:@11028.4]
  wire  storesToCheck_13_3; // @[LoadQueue.scala 131:10:@11029.4]
  wire  _T_10902; // @[LoadQueue.scala 131:81:@11032.4]
  wire  _T_10903; // @[LoadQueue.scala 131:72:@11033.4]
  wire  _T_10905; // @[LoadQueue.scala 132:33:@11034.4]
  wire  _T_10908; // @[LoadQueue.scala 132:41:@11036.4]
  wire  _T_10910; // @[LoadQueue.scala 132:9:@11037.4]
  wire  storesToCheck_13_4; // @[LoadQueue.scala 131:10:@11038.4]
  wire  _T_10916; // @[LoadQueue.scala 131:81:@11041.4]
  wire  _T_10917; // @[LoadQueue.scala 131:72:@11042.4]
  wire  _T_10919; // @[LoadQueue.scala 132:33:@11043.4]
  wire  _T_10922; // @[LoadQueue.scala 132:41:@11045.4]
  wire  _T_10924; // @[LoadQueue.scala 132:9:@11046.4]
  wire  storesToCheck_13_5; // @[LoadQueue.scala 131:10:@11047.4]
  wire  _T_10930; // @[LoadQueue.scala 131:81:@11050.4]
  wire  _T_10931; // @[LoadQueue.scala 131:72:@11051.4]
  wire  _T_10933; // @[LoadQueue.scala 132:33:@11052.4]
  wire  _T_10936; // @[LoadQueue.scala 132:41:@11054.4]
  wire  _T_10938; // @[LoadQueue.scala 132:9:@11055.4]
  wire  storesToCheck_13_6; // @[LoadQueue.scala 131:10:@11056.4]
  wire  _T_10944; // @[LoadQueue.scala 131:81:@11059.4]
  wire  _T_10945; // @[LoadQueue.scala 131:72:@11060.4]
  wire  _T_10947; // @[LoadQueue.scala 132:33:@11061.4]
  wire  _T_10950; // @[LoadQueue.scala 132:41:@11063.4]
  wire  _T_10952; // @[LoadQueue.scala 132:9:@11064.4]
  wire  storesToCheck_13_7; // @[LoadQueue.scala 131:10:@11065.4]
  wire  _T_10958; // @[LoadQueue.scala 131:81:@11068.4]
  wire  _T_10959; // @[LoadQueue.scala 131:72:@11069.4]
  wire  _T_10961; // @[LoadQueue.scala 132:33:@11070.4]
  wire  _T_10964; // @[LoadQueue.scala 132:41:@11072.4]
  wire  _T_10966; // @[LoadQueue.scala 132:9:@11073.4]
  wire  storesToCheck_13_8; // @[LoadQueue.scala 131:10:@11074.4]
  wire  _T_10972; // @[LoadQueue.scala 131:81:@11077.4]
  wire  _T_10973; // @[LoadQueue.scala 131:72:@11078.4]
  wire  _T_10975; // @[LoadQueue.scala 132:33:@11079.4]
  wire  _T_10978; // @[LoadQueue.scala 132:41:@11081.4]
  wire  _T_10980; // @[LoadQueue.scala 132:9:@11082.4]
  wire  storesToCheck_13_9; // @[LoadQueue.scala 131:10:@11083.4]
  wire  _T_10986; // @[LoadQueue.scala 131:81:@11086.4]
  wire  _T_10987; // @[LoadQueue.scala 131:72:@11087.4]
  wire  _T_10989; // @[LoadQueue.scala 132:33:@11088.4]
  wire  _T_10992; // @[LoadQueue.scala 132:41:@11090.4]
  wire  _T_10994; // @[LoadQueue.scala 132:9:@11091.4]
  wire  storesToCheck_13_10; // @[LoadQueue.scala 131:10:@11092.4]
  wire  _T_11000; // @[LoadQueue.scala 131:81:@11095.4]
  wire  _T_11001; // @[LoadQueue.scala 131:72:@11096.4]
  wire  _T_11003; // @[LoadQueue.scala 132:33:@11097.4]
  wire  _T_11006; // @[LoadQueue.scala 132:41:@11099.4]
  wire  _T_11008; // @[LoadQueue.scala 132:9:@11100.4]
  wire  storesToCheck_13_11; // @[LoadQueue.scala 131:10:@11101.4]
  wire  _T_11014; // @[LoadQueue.scala 131:81:@11104.4]
  wire  _T_11015; // @[LoadQueue.scala 131:72:@11105.4]
  wire  _T_11017; // @[LoadQueue.scala 132:33:@11106.4]
  wire  _T_11020; // @[LoadQueue.scala 132:41:@11108.4]
  wire  _T_11022; // @[LoadQueue.scala 132:9:@11109.4]
  wire  storesToCheck_13_12; // @[LoadQueue.scala 131:10:@11110.4]
  wire  _T_11028; // @[LoadQueue.scala 131:81:@11113.4]
  wire  _T_11029; // @[LoadQueue.scala 131:72:@11114.4]
  wire  _T_11031; // @[LoadQueue.scala 132:33:@11115.4]
  wire  _T_11034; // @[LoadQueue.scala 132:41:@11117.4]
  wire  _T_11036; // @[LoadQueue.scala 132:9:@11118.4]
  wire  storesToCheck_13_13; // @[LoadQueue.scala 131:10:@11119.4]
  wire  _T_11042; // @[LoadQueue.scala 131:81:@11122.4]
  wire  _T_11043; // @[LoadQueue.scala 131:72:@11123.4]
  wire  _T_11045; // @[LoadQueue.scala 132:33:@11124.4]
  wire  _T_11048; // @[LoadQueue.scala 132:41:@11126.4]
  wire  _T_11050; // @[LoadQueue.scala 132:9:@11127.4]
  wire  storesToCheck_13_14; // @[LoadQueue.scala 131:10:@11128.4]
  wire  _T_11056; // @[LoadQueue.scala 131:81:@11131.4]
  wire  storesToCheck_13_15; // @[LoadQueue.scala 131:10:@11137.4]
  wire  storesToCheck_14_0; // @[LoadQueue.scala 131:10:@11179.4]
  wire  _T_11106; // @[LoadQueue.scala 131:81:@11182.4]
  wire  _T_11107; // @[LoadQueue.scala 131:72:@11183.4]
  wire  _T_11109; // @[LoadQueue.scala 132:33:@11184.4]
  wire  _T_11112; // @[LoadQueue.scala 132:41:@11186.4]
  wire  _T_11114; // @[LoadQueue.scala 132:9:@11187.4]
  wire  storesToCheck_14_1; // @[LoadQueue.scala 131:10:@11188.4]
  wire  _T_11120; // @[LoadQueue.scala 131:81:@11191.4]
  wire  _T_11121; // @[LoadQueue.scala 131:72:@11192.4]
  wire  _T_11123; // @[LoadQueue.scala 132:33:@11193.4]
  wire  _T_11126; // @[LoadQueue.scala 132:41:@11195.4]
  wire  _T_11128; // @[LoadQueue.scala 132:9:@11196.4]
  wire  storesToCheck_14_2; // @[LoadQueue.scala 131:10:@11197.4]
  wire  _T_11134; // @[LoadQueue.scala 131:81:@11200.4]
  wire  _T_11135; // @[LoadQueue.scala 131:72:@11201.4]
  wire  _T_11137; // @[LoadQueue.scala 132:33:@11202.4]
  wire  _T_11140; // @[LoadQueue.scala 132:41:@11204.4]
  wire  _T_11142; // @[LoadQueue.scala 132:9:@11205.4]
  wire  storesToCheck_14_3; // @[LoadQueue.scala 131:10:@11206.4]
  wire  _T_11148; // @[LoadQueue.scala 131:81:@11209.4]
  wire  _T_11149; // @[LoadQueue.scala 131:72:@11210.4]
  wire  _T_11151; // @[LoadQueue.scala 132:33:@11211.4]
  wire  _T_11154; // @[LoadQueue.scala 132:41:@11213.4]
  wire  _T_11156; // @[LoadQueue.scala 132:9:@11214.4]
  wire  storesToCheck_14_4; // @[LoadQueue.scala 131:10:@11215.4]
  wire  _T_11162; // @[LoadQueue.scala 131:81:@11218.4]
  wire  _T_11163; // @[LoadQueue.scala 131:72:@11219.4]
  wire  _T_11165; // @[LoadQueue.scala 132:33:@11220.4]
  wire  _T_11168; // @[LoadQueue.scala 132:41:@11222.4]
  wire  _T_11170; // @[LoadQueue.scala 132:9:@11223.4]
  wire  storesToCheck_14_5; // @[LoadQueue.scala 131:10:@11224.4]
  wire  _T_11176; // @[LoadQueue.scala 131:81:@11227.4]
  wire  _T_11177; // @[LoadQueue.scala 131:72:@11228.4]
  wire  _T_11179; // @[LoadQueue.scala 132:33:@11229.4]
  wire  _T_11182; // @[LoadQueue.scala 132:41:@11231.4]
  wire  _T_11184; // @[LoadQueue.scala 132:9:@11232.4]
  wire  storesToCheck_14_6; // @[LoadQueue.scala 131:10:@11233.4]
  wire  _T_11190; // @[LoadQueue.scala 131:81:@11236.4]
  wire  _T_11191; // @[LoadQueue.scala 131:72:@11237.4]
  wire  _T_11193; // @[LoadQueue.scala 132:33:@11238.4]
  wire  _T_11196; // @[LoadQueue.scala 132:41:@11240.4]
  wire  _T_11198; // @[LoadQueue.scala 132:9:@11241.4]
  wire  storesToCheck_14_7; // @[LoadQueue.scala 131:10:@11242.4]
  wire  _T_11204; // @[LoadQueue.scala 131:81:@11245.4]
  wire  _T_11205; // @[LoadQueue.scala 131:72:@11246.4]
  wire  _T_11207; // @[LoadQueue.scala 132:33:@11247.4]
  wire  _T_11210; // @[LoadQueue.scala 132:41:@11249.4]
  wire  _T_11212; // @[LoadQueue.scala 132:9:@11250.4]
  wire  storesToCheck_14_8; // @[LoadQueue.scala 131:10:@11251.4]
  wire  _T_11218; // @[LoadQueue.scala 131:81:@11254.4]
  wire  _T_11219; // @[LoadQueue.scala 131:72:@11255.4]
  wire  _T_11221; // @[LoadQueue.scala 132:33:@11256.4]
  wire  _T_11224; // @[LoadQueue.scala 132:41:@11258.4]
  wire  _T_11226; // @[LoadQueue.scala 132:9:@11259.4]
  wire  storesToCheck_14_9; // @[LoadQueue.scala 131:10:@11260.4]
  wire  _T_11232; // @[LoadQueue.scala 131:81:@11263.4]
  wire  _T_11233; // @[LoadQueue.scala 131:72:@11264.4]
  wire  _T_11235; // @[LoadQueue.scala 132:33:@11265.4]
  wire  _T_11238; // @[LoadQueue.scala 132:41:@11267.4]
  wire  _T_11240; // @[LoadQueue.scala 132:9:@11268.4]
  wire  storesToCheck_14_10; // @[LoadQueue.scala 131:10:@11269.4]
  wire  _T_11246; // @[LoadQueue.scala 131:81:@11272.4]
  wire  _T_11247; // @[LoadQueue.scala 131:72:@11273.4]
  wire  _T_11249; // @[LoadQueue.scala 132:33:@11274.4]
  wire  _T_11252; // @[LoadQueue.scala 132:41:@11276.4]
  wire  _T_11254; // @[LoadQueue.scala 132:9:@11277.4]
  wire  storesToCheck_14_11; // @[LoadQueue.scala 131:10:@11278.4]
  wire  _T_11260; // @[LoadQueue.scala 131:81:@11281.4]
  wire  _T_11261; // @[LoadQueue.scala 131:72:@11282.4]
  wire  _T_11263; // @[LoadQueue.scala 132:33:@11283.4]
  wire  _T_11266; // @[LoadQueue.scala 132:41:@11285.4]
  wire  _T_11268; // @[LoadQueue.scala 132:9:@11286.4]
  wire  storesToCheck_14_12; // @[LoadQueue.scala 131:10:@11287.4]
  wire  _T_11274; // @[LoadQueue.scala 131:81:@11290.4]
  wire  _T_11275; // @[LoadQueue.scala 131:72:@11291.4]
  wire  _T_11277; // @[LoadQueue.scala 132:33:@11292.4]
  wire  _T_11280; // @[LoadQueue.scala 132:41:@11294.4]
  wire  _T_11282; // @[LoadQueue.scala 132:9:@11295.4]
  wire  storesToCheck_14_13; // @[LoadQueue.scala 131:10:@11296.4]
  wire  _T_11288; // @[LoadQueue.scala 131:81:@11299.4]
  wire  _T_11289; // @[LoadQueue.scala 131:72:@11300.4]
  wire  _T_11291; // @[LoadQueue.scala 132:33:@11301.4]
  wire  _T_11294; // @[LoadQueue.scala 132:41:@11303.4]
  wire  _T_11296; // @[LoadQueue.scala 132:9:@11304.4]
  wire  storesToCheck_14_14; // @[LoadQueue.scala 131:10:@11305.4]
  wire  _T_11302; // @[LoadQueue.scala 131:81:@11308.4]
  wire  storesToCheck_14_15; // @[LoadQueue.scala 131:10:@11314.4]
  wire  storesToCheck_15_0; // @[LoadQueue.scala 131:10:@11356.4]
  wire  _T_11352; // @[LoadQueue.scala 131:81:@11359.4]
  wire  _T_11353; // @[LoadQueue.scala 131:72:@11360.4]
  wire  _T_11355; // @[LoadQueue.scala 132:33:@11361.4]
  wire  _T_11358; // @[LoadQueue.scala 132:41:@11363.4]
  wire  _T_11360; // @[LoadQueue.scala 132:9:@11364.4]
  wire  storesToCheck_15_1; // @[LoadQueue.scala 131:10:@11365.4]
  wire  _T_11366; // @[LoadQueue.scala 131:81:@11368.4]
  wire  _T_11367; // @[LoadQueue.scala 131:72:@11369.4]
  wire  _T_11369; // @[LoadQueue.scala 132:33:@11370.4]
  wire  _T_11372; // @[LoadQueue.scala 132:41:@11372.4]
  wire  _T_11374; // @[LoadQueue.scala 132:9:@11373.4]
  wire  storesToCheck_15_2; // @[LoadQueue.scala 131:10:@11374.4]
  wire  _T_11380; // @[LoadQueue.scala 131:81:@11377.4]
  wire  _T_11381; // @[LoadQueue.scala 131:72:@11378.4]
  wire  _T_11383; // @[LoadQueue.scala 132:33:@11379.4]
  wire  _T_11386; // @[LoadQueue.scala 132:41:@11381.4]
  wire  _T_11388; // @[LoadQueue.scala 132:9:@11382.4]
  wire  storesToCheck_15_3; // @[LoadQueue.scala 131:10:@11383.4]
  wire  _T_11394; // @[LoadQueue.scala 131:81:@11386.4]
  wire  _T_11395; // @[LoadQueue.scala 131:72:@11387.4]
  wire  _T_11397; // @[LoadQueue.scala 132:33:@11388.4]
  wire  _T_11400; // @[LoadQueue.scala 132:41:@11390.4]
  wire  _T_11402; // @[LoadQueue.scala 132:9:@11391.4]
  wire  storesToCheck_15_4; // @[LoadQueue.scala 131:10:@11392.4]
  wire  _T_11408; // @[LoadQueue.scala 131:81:@11395.4]
  wire  _T_11409; // @[LoadQueue.scala 131:72:@11396.4]
  wire  _T_11411; // @[LoadQueue.scala 132:33:@11397.4]
  wire  _T_11414; // @[LoadQueue.scala 132:41:@11399.4]
  wire  _T_11416; // @[LoadQueue.scala 132:9:@11400.4]
  wire  storesToCheck_15_5; // @[LoadQueue.scala 131:10:@11401.4]
  wire  _T_11422; // @[LoadQueue.scala 131:81:@11404.4]
  wire  _T_11423; // @[LoadQueue.scala 131:72:@11405.4]
  wire  _T_11425; // @[LoadQueue.scala 132:33:@11406.4]
  wire  _T_11428; // @[LoadQueue.scala 132:41:@11408.4]
  wire  _T_11430; // @[LoadQueue.scala 132:9:@11409.4]
  wire  storesToCheck_15_6; // @[LoadQueue.scala 131:10:@11410.4]
  wire  _T_11436; // @[LoadQueue.scala 131:81:@11413.4]
  wire  _T_11437; // @[LoadQueue.scala 131:72:@11414.4]
  wire  _T_11439; // @[LoadQueue.scala 132:33:@11415.4]
  wire  _T_11442; // @[LoadQueue.scala 132:41:@11417.4]
  wire  _T_11444; // @[LoadQueue.scala 132:9:@11418.4]
  wire  storesToCheck_15_7; // @[LoadQueue.scala 131:10:@11419.4]
  wire  _T_11450; // @[LoadQueue.scala 131:81:@11422.4]
  wire  _T_11451; // @[LoadQueue.scala 131:72:@11423.4]
  wire  _T_11453; // @[LoadQueue.scala 132:33:@11424.4]
  wire  _T_11456; // @[LoadQueue.scala 132:41:@11426.4]
  wire  _T_11458; // @[LoadQueue.scala 132:9:@11427.4]
  wire  storesToCheck_15_8; // @[LoadQueue.scala 131:10:@11428.4]
  wire  _T_11464; // @[LoadQueue.scala 131:81:@11431.4]
  wire  _T_11465; // @[LoadQueue.scala 131:72:@11432.4]
  wire  _T_11467; // @[LoadQueue.scala 132:33:@11433.4]
  wire  _T_11470; // @[LoadQueue.scala 132:41:@11435.4]
  wire  _T_11472; // @[LoadQueue.scala 132:9:@11436.4]
  wire  storesToCheck_15_9; // @[LoadQueue.scala 131:10:@11437.4]
  wire  _T_11478; // @[LoadQueue.scala 131:81:@11440.4]
  wire  _T_11479; // @[LoadQueue.scala 131:72:@11441.4]
  wire  _T_11481; // @[LoadQueue.scala 132:33:@11442.4]
  wire  _T_11484; // @[LoadQueue.scala 132:41:@11444.4]
  wire  _T_11486; // @[LoadQueue.scala 132:9:@11445.4]
  wire  storesToCheck_15_10; // @[LoadQueue.scala 131:10:@11446.4]
  wire  _T_11492; // @[LoadQueue.scala 131:81:@11449.4]
  wire  _T_11493; // @[LoadQueue.scala 131:72:@11450.4]
  wire  _T_11495; // @[LoadQueue.scala 132:33:@11451.4]
  wire  _T_11498; // @[LoadQueue.scala 132:41:@11453.4]
  wire  _T_11500; // @[LoadQueue.scala 132:9:@11454.4]
  wire  storesToCheck_15_11; // @[LoadQueue.scala 131:10:@11455.4]
  wire  _T_11506; // @[LoadQueue.scala 131:81:@11458.4]
  wire  _T_11507; // @[LoadQueue.scala 131:72:@11459.4]
  wire  _T_11509; // @[LoadQueue.scala 132:33:@11460.4]
  wire  _T_11512; // @[LoadQueue.scala 132:41:@11462.4]
  wire  _T_11514; // @[LoadQueue.scala 132:9:@11463.4]
  wire  storesToCheck_15_12; // @[LoadQueue.scala 131:10:@11464.4]
  wire  _T_11520; // @[LoadQueue.scala 131:81:@11467.4]
  wire  _T_11521; // @[LoadQueue.scala 131:72:@11468.4]
  wire  _T_11523; // @[LoadQueue.scala 132:33:@11469.4]
  wire  _T_11526; // @[LoadQueue.scala 132:41:@11471.4]
  wire  _T_11528; // @[LoadQueue.scala 132:9:@11472.4]
  wire  storesToCheck_15_13; // @[LoadQueue.scala 131:10:@11473.4]
  wire  _T_11534; // @[LoadQueue.scala 131:81:@11476.4]
  wire  _T_11535; // @[LoadQueue.scala 131:72:@11477.4]
  wire  _T_11537; // @[LoadQueue.scala 132:33:@11478.4]
  wire  _T_11540; // @[LoadQueue.scala 132:41:@11480.4]
  wire  _T_11542; // @[LoadQueue.scala 132:9:@11481.4]
  wire  storesToCheck_15_14; // @[LoadQueue.scala 131:10:@11482.4]
  wire  _T_11548; // @[LoadQueue.scala 131:81:@11485.4]
  wire  storesToCheck_15_15; // @[LoadQueue.scala 131:10:@11491.4]
  wire  _T_12810; // @[LoadQueue.scala 141:18:@11526.4]
  wire  entriesToCheck_0_0; // @[LoadQueue.scala 141:26:@11527.4]
  wire  _T_12812; // @[LoadQueue.scala 141:18:@11528.4]
  wire  entriesToCheck_0_1; // @[LoadQueue.scala 141:26:@11529.4]
  wire  _T_12814; // @[LoadQueue.scala 141:18:@11530.4]
  wire  entriesToCheck_0_2; // @[LoadQueue.scala 141:26:@11531.4]
  wire  _T_12816; // @[LoadQueue.scala 141:18:@11532.4]
  wire  entriesToCheck_0_3; // @[LoadQueue.scala 141:26:@11533.4]
  wire  _T_12818; // @[LoadQueue.scala 141:18:@11534.4]
  wire  entriesToCheck_0_4; // @[LoadQueue.scala 141:26:@11535.4]
  wire  _T_12820; // @[LoadQueue.scala 141:18:@11536.4]
  wire  entriesToCheck_0_5; // @[LoadQueue.scala 141:26:@11537.4]
  wire  _T_12822; // @[LoadQueue.scala 141:18:@11538.4]
  wire  entriesToCheck_0_6; // @[LoadQueue.scala 141:26:@11539.4]
  wire  _T_12824; // @[LoadQueue.scala 141:18:@11540.4]
  wire  entriesToCheck_0_7; // @[LoadQueue.scala 141:26:@11541.4]
  wire  _T_12826; // @[LoadQueue.scala 141:18:@11542.4]
  wire  entriesToCheck_0_8; // @[LoadQueue.scala 141:26:@11543.4]
  wire  _T_12828; // @[LoadQueue.scala 141:18:@11544.4]
  wire  entriesToCheck_0_9; // @[LoadQueue.scala 141:26:@11545.4]
  wire  _T_12830; // @[LoadQueue.scala 141:18:@11546.4]
  wire  entriesToCheck_0_10; // @[LoadQueue.scala 141:26:@11547.4]
  wire  _T_12832; // @[LoadQueue.scala 141:18:@11548.4]
  wire  entriesToCheck_0_11; // @[LoadQueue.scala 141:26:@11549.4]
  wire  _T_12834; // @[LoadQueue.scala 141:18:@11550.4]
  wire  entriesToCheck_0_12; // @[LoadQueue.scala 141:26:@11551.4]
  wire  _T_12836; // @[LoadQueue.scala 141:18:@11552.4]
  wire  entriesToCheck_0_13; // @[LoadQueue.scala 141:26:@11553.4]
  wire  _T_12838; // @[LoadQueue.scala 141:18:@11554.4]
  wire  entriesToCheck_0_14; // @[LoadQueue.scala 141:26:@11555.4]
  wire  _T_12840; // @[LoadQueue.scala 141:18:@11556.4]
  wire  entriesToCheck_0_15; // @[LoadQueue.scala 141:26:@11557.4]
  wire  _T_12842; // @[LoadQueue.scala 141:18:@11574.4]
  wire  entriesToCheck_1_0; // @[LoadQueue.scala 141:26:@11575.4]
  wire  _T_12844; // @[LoadQueue.scala 141:18:@11576.4]
  wire  entriesToCheck_1_1; // @[LoadQueue.scala 141:26:@11577.4]
  wire  _T_12846; // @[LoadQueue.scala 141:18:@11578.4]
  wire  entriesToCheck_1_2; // @[LoadQueue.scala 141:26:@11579.4]
  wire  _T_12848; // @[LoadQueue.scala 141:18:@11580.4]
  wire  entriesToCheck_1_3; // @[LoadQueue.scala 141:26:@11581.4]
  wire  _T_12850; // @[LoadQueue.scala 141:18:@11582.4]
  wire  entriesToCheck_1_4; // @[LoadQueue.scala 141:26:@11583.4]
  wire  _T_12852; // @[LoadQueue.scala 141:18:@11584.4]
  wire  entriesToCheck_1_5; // @[LoadQueue.scala 141:26:@11585.4]
  wire  _T_12854; // @[LoadQueue.scala 141:18:@11586.4]
  wire  entriesToCheck_1_6; // @[LoadQueue.scala 141:26:@11587.4]
  wire  _T_12856; // @[LoadQueue.scala 141:18:@11588.4]
  wire  entriesToCheck_1_7; // @[LoadQueue.scala 141:26:@11589.4]
  wire  _T_12858; // @[LoadQueue.scala 141:18:@11590.4]
  wire  entriesToCheck_1_8; // @[LoadQueue.scala 141:26:@11591.4]
  wire  _T_12860; // @[LoadQueue.scala 141:18:@11592.4]
  wire  entriesToCheck_1_9; // @[LoadQueue.scala 141:26:@11593.4]
  wire  _T_12862; // @[LoadQueue.scala 141:18:@11594.4]
  wire  entriesToCheck_1_10; // @[LoadQueue.scala 141:26:@11595.4]
  wire  _T_12864; // @[LoadQueue.scala 141:18:@11596.4]
  wire  entriesToCheck_1_11; // @[LoadQueue.scala 141:26:@11597.4]
  wire  _T_12866; // @[LoadQueue.scala 141:18:@11598.4]
  wire  entriesToCheck_1_12; // @[LoadQueue.scala 141:26:@11599.4]
  wire  _T_12868; // @[LoadQueue.scala 141:18:@11600.4]
  wire  entriesToCheck_1_13; // @[LoadQueue.scala 141:26:@11601.4]
  wire  _T_12870; // @[LoadQueue.scala 141:18:@11602.4]
  wire  entriesToCheck_1_14; // @[LoadQueue.scala 141:26:@11603.4]
  wire  _T_12872; // @[LoadQueue.scala 141:18:@11604.4]
  wire  entriesToCheck_1_15; // @[LoadQueue.scala 141:26:@11605.4]
  wire  _T_12874; // @[LoadQueue.scala 141:18:@11622.4]
  wire  entriesToCheck_2_0; // @[LoadQueue.scala 141:26:@11623.4]
  wire  _T_12876; // @[LoadQueue.scala 141:18:@11624.4]
  wire  entriesToCheck_2_1; // @[LoadQueue.scala 141:26:@11625.4]
  wire  _T_12878; // @[LoadQueue.scala 141:18:@11626.4]
  wire  entriesToCheck_2_2; // @[LoadQueue.scala 141:26:@11627.4]
  wire  _T_12880; // @[LoadQueue.scala 141:18:@11628.4]
  wire  entriesToCheck_2_3; // @[LoadQueue.scala 141:26:@11629.4]
  wire  _T_12882; // @[LoadQueue.scala 141:18:@11630.4]
  wire  entriesToCheck_2_4; // @[LoadQueue.scala 141:26:@11631.4]
  wire  _T_12884; // @[LoadQueue.scala 141:18:@11632.4]
  wire  entriesToCheck_2_5; // @[LoadQueue.scala 141:26:@11633.4]
  wire  _T_12886; // @[LoadQueue.scala 141:18:@11634.4]
  wire  entriesToCheck_2_6; // @[LoadQueue.scala 141:26:@11635.4]
  wire  _T_12888; // @[LoadQueue.scala 141:18:@11636.4]
  wire  entriesToCheck_2_7; // @[LoadQueue.scala 141:26:@11637.4]
  wire  _T_12890; // @[LoadQueue.scala 141:18:@11638.4]
  wire  entriesToCheck_2_8; // @[LoadQueue.scala 141:26:@11639.4]
  wire  _T_12892; // @[LoadQueue.scala 141:18:@11640.4]
  wire  entriesToCheck_2_9; // @[LoadQueue.scala 141:26:@11641.4]
  wire  _T_12894; // @[LoadQueue.scala 141:18:@11642.4]
  wire  entriesToCheck_2_10; // @[LoadQueue.scala 141:26:@11643.4]
  wire  _T_12896; // @[LoadQueue.scala 141:18:@11644.4]
  wire  entriesToCheck_2_11; // @[LoadQueue.scala 141:26:@11645.4]
  wire  _T_12898; // @[LoadQueue.scala 141:18:@11646.4]
  wire  entriesToCheck_2_12; // @[LoadQueue.scala 141:26:@11647.4]
  wire  _T_12900; // @[LoadQueue.scala 141:18:@11648.4]
  wire  entriesToCheck_2_13; // @[LoadQueue.scala 141:26:@11649.4]
  wire  _T_12902; // @[LoadQueue.scala 141:18:@11650.4]
  wire  entriesToCheck_2_14; // @[LoadQueue.scala 141:26:@11651.4]
  wire  _T_12904; // @[LoadQueue.scala 141:18:@11652.4]
  wire  entriesToCheck_2_15; // @[LoadQueue.scala 141:26:@11653.4]
  wire  _T_12906; // @[LoadQueue.scala 141:18:@11670.4]
  wire  entriesToCheck_3_0; // @[LoadQueue.scala 141:26:@11671.4]
  wire  _T_12908; // @[LoadQueue.scala 141:18:@11672.4]
  wire  entriesToCheck_3_1; // @[LoadQueue.scala 141:26:@11673.4]
  wire  _T_12910; // @[LoadQueue.scala 141:18:@11674.4]
  wire  entriesToCheck_3_2; // @[LoadQueue.scala 141:26:@11675.4]
  wire  _T_12912; // @[LoadQueue.scala 141:18:@11676.4]
  wire  entriesToCheck_3_3; // @[LoadQueue.scala 141:26:@11677.4]
  wire  _T_12914; // @[LoadQueue.scala 141:18:@11678.4]
  wire  entriesToCheck_3_4; // @[LoadQueue.scala 141:26:@11679.4]
  wire  _T_12916; // @[LoadQueue.scala 141:18:@11680.4]
  wire  entriesToCheck_3_5; // @[LoadQueue.scala 141:26:@11681.4]
  wire  _T_12918; // @[LoadQueue.scala 141:18:@11682.4]
  wire  entriesToCheck_3_6; // @[LoadQueue.scala 141:26:@11683.4]
  wire  _T_12920; // @[LoadQueue.scala 141:18:@11684.4]
  wire  entriesToCheck_3_7; // @[LoadQueue.scala 141:26:@11685.4]
  wire  _T_12922; // @[LoadQueue.scala 141:18:@11686.4]
  wire  entriesToCheck_3_8; // @[LoadQueue.scala 141:26:@11687.4]
  wire  _T_12924; // @[LoadQueue.scala 141:18:@11688.4]
  wire  entriesToCheck_3_9; // @[LoadQueue.scala 141:26:@11689.4]
  wire  _T_12926; // @[LoadQueue.scala 141:18:@11690.4]
  wire  entriesToCheck_3_10; // @[LoadQueue.scala 141:26:@11691.4]
  wire  _T_12928; // @[LoadQueue.scala 141:18:@11692.4]
  wire  entriesToCheck_3_11; // @[LoadQueue.scala 141:26:@11693.4]
  wire  _T_12930; // @[LoadQueue.scala 141:18:@11694.4]
  wire  entriesToCheck_3_12; // @[LoadQueue.scala 141:26:@11695.4]
  wire  _T_12932; // @[LoadQueue.scala 141:18:@11696.4]
  wire  entriesToCheck_3_13; // @[LoadQueue.scala 141:26:@11697.4]
  wire  _T_12934; // @[LoadQueue.scala 141:18:@11698.4]
  wire  entriesToCheck_3_14; // @[LoadQueue.scala 141:26:@11699.4]
  wire  _T_12936; // @[LoadQueue.scala 141:18:@11700.4]
  wire  entriesToCheck_3_15; // @[LoadQueue.scala 141:26:@11701.4]
  wire  _T_12938; // @[LoadQueue.scala 141:18:@11718.4]
  wire  entriesToCheck_4_0; // @[LoadQueue.scala 141:26:@11719.4]
  wire  _T_12940; // @[LoadQueue.scala 141:18:@11720.4]
  wire  entriesToCheck_4_1; // @[LoadQueue.scala 141:26:@11721.4]
  wire  _T_12942; // @[LoadQueue.scala 141:18:@11722.4]
  wire  entriesToCheck_4_2; // @[LoadQueue.scala 141:26:@11723.4]
  wire  _T_12944; // @[LoadQueue.scala 141:18:@11724.4]
  wire  entriesToCheck_4_3; // @[LoadQueue.scala 141:26:@11725.4]
  wire  _T_12946; // @[LoadQueue.scala 141:18:@11726.4]
  wire  entriesToCheck_4_4; // @[LoadQueue.scala 141:26:@11727.4]
  wire  _T_12948; // @[LoadQueue.scala 141:18:@11728.4]
  wire  entriesToCheck_4_5; // @[LoadQueue.scala 141:26:@11729.4]
  wire  _T_12950; // @[LoadQueue.scala 141:18:@11730.4]
  wire  entriesToCheck_4_6; // @[LoadQueue.scala 141:26:@11731.4]
  wire  _T_12952; // @[LoadQueue.scala 141:18:@11732.4]
  wire  entriesToCheck_4_7; // @[LoadQueue.scala 141:26:@11733.4]
  wire  _T_12954; // @[LoadQueue.scala 141:18:@11734.4]
  wire  entriesToCheck_4_8; // @[LoadQueue.scala 141:26:@11735.4]
  wire  _T_12956; // @[LoadQueue.scala 141:18:@11736.4]
  wire  entriesToCheck_4_9; // @[LoadQueue.scala 141:26:@11737.4]
  wire  _T_12958; // @[LoadQueue.scala 141:18:@11738.4]
  wire  entriesToCheck_4_10; // @[LoadQueue.scala 141:26:@11739.4]
  wire  _T_12960; // @[LoadQueue.scala 141:18:@11740.4]
  wire  entriesToCheck_4_11; // @[LoadQueue.scala 141:26:@11741.4]
  wire  _T_12962; // @[LoadQueue.scala 141:18:@11742.4]
  wire  entriesToCheck_4_12; // @[LoadQueue.scala 141:26:@11743.4]
  wire  _T_12964; // @[LoadQueue.scala 141:18:@11744.4]
  wire  entriesToCheck_4_13; // @[LoadQueue.scala 141:26:@11745.4]
  wire  _T_12966; // @[LoadQueue.scala 141:18:@11746.4]
  wire  entriesToCheck_4_14; // @[LoadQueue.scala 141:26:@11747.4]
  wire  _T_12968; // @[LoadQueue.scala 141:18:@11748.4]
  wire  entriesToCheck_4_15; // @[LoadQueue.scala 141:26:@11749.4]
  wire  _T_12970; // @[LoadQueue.scala 141:18:@11766.4]
  wire  entriesToCheck_5_0; // @[LoadQueue.scala 141:26:@11767.4]
  wire  _T_12972; // @[LoadQueue.scala 141:18:@11768.4]
  wire  entriesToCheck_5_1; // @[LoadQueue.scala 141:26:@11769.4]
  wire  _T_12974; // @[LoadQueue.scala 141:18:@11770.4]
  wire  entriesToCheck_5_2; // @[LoadQueue.scala 141:26:@11771.4]
  wire  _T_12976; // @[LoadQueue.scala 141:18:@11772.4]
  wire  entriesToCheck_5_3; // @[LoadQueue.scala 141:26:@11773.4]
  wire  _T_12978; // @[LoadQueue.scala 141:18:@11774.4]
  wire  entriesToCheck_5_4; // @[LoadQueue.scala 141:26:@11775.4]
  wire  _T_12980; // @[LoadQueue.scala 141:18:@11776.4]
  wire  entriesToCheck_5_5; // @[LoadQueue.scala 141:26:@11777.4]
  wire  _T_12982; // @[LoadQueue.scala 141:18:@11778.4]
  wire  entriesToCheck_5_6; // @[LoadQueue.scala 141:26:@11779.4]
  wire  _T_12984; // @[LoadQueue.scala 141:18:@11780.4]
  wire  entriesToCheck_5_7; // @[LoadQueue.scala 141:26:@11781.4]
  wire  _T_12986; // @[LoadQueue.scala 141:18:@11782.4]
  wire  entriesToCheck_5_8; // @[LoadQueue.scala 141:26:@11783.4]
  wire  _T_12988; // @[LoadQueue.scala 141:18:@11784.4]
  wire  entriesToCheck_5_9; // @[LoadQueue.scala 141:26:@11785.4]
  wire  _T_12990; // @[LoadQueue.scala 141:18:@11786.4]
  wire  entriesToCheck_5_10; // @[LoadQueue.scala 141:26:@11787.4]
  wire  _T_12992; // @[LoadQueue.scala 141:18:@11788.4]
  wire  entriesToCheck_5_11; // @[LoadQueue.scala 141:26:@11789.4]
  wire  _T_12994; // @[LoadQueue.scala 141:18:@11790.4]
  wire  entriesToCheck_5_12; // @[LoadQueue.scala 141:26:@11791.4]
  wire  _T_12996; // @[LoadQueue.scala 141:18:@11792.4]
  wire  entriesToCheck_5_13; // @[LoadQueue.scala 141:26:@11793.4]
  wire  _T_12998; // @[LoadQueue.scala 141:18:@11794.4]
  wire  entriesToCheck_5_14; // @[LoadQueue.scala 141:26:@11795.4]
  wire  _T_13000; // @[LoadQueue.scala 141:18:@11796.4]
  wire  entriesToCheck_5_15; // @[LoadQueue.scala 141:26:@11797.4]
  wire  _T_13002; // @[LoadQueue.scala 141:18:@11814.4]
  wire  entriesToCheck_6_0; // @[LoadQueue.scala 141:26:@11815.4]
  wire  _T_13004; // @[LoadQueue.scala 141:18:@11816.4]
  wire  entriesToCheck_6_1; // @[LoadQueue.scala 141:26:@11817.4]
  wire  _T_13006; // @[LoadQueue.scala 141:18:@11818.4]
  wire  entriesToCheck_6_2; // @[LoadQueue.scala 141:26:@11819.4]
  wire  _T_13008; // @[LoadQueue.scala 141:18:@11820.4]
  wire  entriesToCheck_6_3; // @[LoadQueue.scala 141:26:@11821.4]
  wire  _T_13010; // @[LoadQueue.scala 141:18:@11822.4]
  wire  entriesToCheck_6_4; // @[LoadQueue.scala 141:26:@11823.4]
  wire  _T_13012; // @[LoadQueue.scala 141:18:@11824.4]
  wire  entriesToCheck_6_5; // @[LoadQueue.scala 141:26:@11825.4]
  wire  _T_13014; // @[LoadQueue.scala 141:18:@11826.4]
  wire  entriesToCheck_6_6; // @[LoadQueue.scala 141:26:@11827.4]
  wire  _T_13016; // @[LoadQueue.scala 141:18:@11828.4]
  wire  entriesToCheck_6_7; // @[LoadQueue.scala 141:26:@11829.4]
  wire  _T_13018; // @[LoadQueue.scala 141:18:@11830.4]
  wire  entriesToCheck_6_8; // @[LoadQueue.scala 141:26:@11831.4]
  wire  _T_13020; // @[LoadQueue.scala 141:18:@11832.4]
  wire  entriesToCheck_6_9; // @[LoadQueue.scala 141:26:@11833.4]
  wire  _T_13022; // @[LoadQueue.scala 141:18:@11834.4]
  wire  entriesToCheck_6_10; // @[LoadQueue.scala 141:26:@11835.4]
  wire  _T_13024; // @[LoadQueue.scala 141:18:@11836.4]
  wire  entriesToCheck_6_11; // @[LoadQueue.scala 141:26:@11837.4]
  wire  _T_13026; // @[LoadQueue.scala 141:18:@11838.4]
  wire  entriesToCheck_6_12; // @[LoadQueue.scala 141:26:@11839.4]
  wire  _T_13028; // @[LoadQueue.scala 141:18:@11840.4]
  wire  entriesToCheck_6_13; // @[LoadQueue.scala 141:26:@11841.4]
  wire  _T_13030; // @[LoadQueue.scala 141:18:@11842.4]
  wire  entriesToCheck_6_14; // @[LoadQueue.scala 141:26:@11843.4]
  wire  _T_13032; // @[LoadQueue.scala 141:18:@11844.4]
  wire  entriesToCheck_6_15; // @[LoadQueue.scala 141:26:@11845.4]
  wire  _T_13034; // @[LoadQueue.scala 141:18:@11862.4]
  wire  entriesToCheck_7_0; // @[LoadQueue.scala 141:26:@11863.4]
  wire  _T_13036; // @[LoadQueue.scala 141:18:@11864.4]
  wire  entriesToCheck_7_1; // @[LoadQueue.scala 141:26:@11865.4]
  wire  _T_13038; // @[LoadQueue.scala 141:18:@11866.4]
  wire  entriesToCheck_7_2; // @[LoadQueue.scala 141:26:@11867.4]
  wire  _T_13040; // @[LoadQueue.scala 141:18:@11868.4]
  wire  entriesToCheck_7_3; // @[LoadQueue.scala 141:26:@11869.4]
  wire  _T_13042; // @[LoadQueue.scala 141:18:@11870.4]
  wire  entriesToCheck_7_4; // @[LoadQueue.scala 141:26:@11871.4]
  wire  _T_13044; // @[LoadQueue.scala 141:18:@11872.4]
  wire  entriesToCheck_7_5; // @[LoadQueue.scala 141:26:@11873.4]
  wire  _T_13046; // @[LoadQueue.scala 141:18:@11874.4]
  wire  entriesToCheck_7_6; // @[LoadQueue.scala 141:26:@11875.4]
  wire  _T_13048; // @[LoadQueue.scala 141:18:@11876.4]
  wire  entriesToCheck_7_7; // @[LoadQueue.scala 141:26:@11877.4]
  wire  _T_13050; // @[LoadQueue.scala 141:18:@11878.4]
  wire  entriesToCheck_7_8; // @[LoadQueue.scala 141:26:@11879.4]
  wire  _T_13052; // @[LoadQueue.scala 141:18:@11880.4]
  wire  entriesToCheck_7_9; // @[LoadQueue.scala 141:26:@11881.4]
  wire  _T_13054; // @[LoadQueue.scala 141:18:@11882.4]
  wire  entriesToCheck_7_10; // @[LoadQueue.scala 141:26:@11883.4]
  wire  _T_13056; // @[LoadQueue.scala 141:18:@11884.4]
  wire  entriesToCheck_7_11; // @[LoadQueue.scala 141:26:@11885.4]
  wire  _T_13058; // @[LoadQueue.scala 141:18:@11886.4]
  wire  entriesToCheck_7_12; // @[LoadQueue.scala 141:26:@11887.4]
  wire  _T_13060; // @[LoadQueue.scala 141:18:@11888.4]
  wire  entriesToCheck_7_13; // @[LoadQueue.scala 141:26:@11889.4]
  wire  _T_13062; // @[LoadQueue.scala 141:18:@11890.4]
  wire  entriesToCheck_7_14; // @[LoadQueue.scala 141:26:@11891.4]
  wire  _T_13064; // @[LoadQueue.scala 141:18:@11892.4]
  wire  entriesToCheck_7_15; // @[LoadQueue.scala 141:26:@11893.4]
  wire  _T_13066; // @[LoadQueue.scala 141:18:@11910.4]
  wire  entriesToCheck_8_0; // @[LoadQueue.scala 141:26:@11911.4]
  wire  _T_13068; // @[LoadQueue.scala 141:18:@11912.4]
  wire  entriesToCheck_8_1; // @[LoadQueue.scala 141:26:@11913.4]
  wire  _T_13070; // @[LoadQueue.scala 141:18:@11914.4]
  wire  entriesToCheck_8_2; // @[LoadQueue.scala 141:26:@11915.4]
  wire  _T_13072; // @[LoadQueue.scala 141:18:@11916.4]
  wire  entriesToCheck_8_3; // @[LoadQueue.scala 141:26:@11917.4]
  wire  _T_13074; // @[LoadQueue.scala 141:18:@11918.4]
  wire  entriesToCheck_8_4; // @[LoadQueue.scala 141:26:@11919.4]
  wire  _T_13076; // @[LoadQueue.scala 141:18:@11920.4]
  wire  entriesToCheck_8_5; // @[LoadQueue.scala 141:26:@11921.4]
  wire  _T_13078; // @[LoadQueue.scala 141:18:@11922.4]
  wire  entriesToCheck_8_6; // @[LoadQueue.scala 141:26:@11923.4]
  wire  _T_13080; // @[LoadQueue.scala 141:18:@11924.4]
  wire  entriesToCheck_8_7; // @[LoadQueue.scala 141:26:@11925.4]
  wire  _T_13082; // @[LoadQueue.scala 141:18:@11926.4]
  wire  entriesToCheck_8_8; // @[LoadQueue.scala 141:26:@11927.4]
  wire  _T_13084; // @[LoadQueue.scala 141:18:@11928.4]
  wire  entriesToCheck_8_9; // @[LoadQueue.scala 141:26:@11929.4]
  wire  _T_13086; // @[LoadQueue.scala 141:18:@11930.4]
  wire  entriesToCheck_8_10; // @[LoadQueue.scala 141:26:@11931.4]
  wire  _T_13088; // @[LoadQueue.scala 141:18:@11932.4]
  wire  entriesToCheck_8_11; // @[LoadQueue.scala 141:26:@11933.4]
  wire  _T_13090; // @[LoadQueue.scala 141:18:@11934.4]
  wire  entriesToCheck_8_12; // @[LoadQueue.scala 141:26:@11935.4]
  wire  _T_13092; // @[LoadQueue.scala 141:18:@11936.4]
  wire  entriesToCheck_8_13; // @[LoadQueue.scala 141:26:@11937.4]
  wire  _T_13094; // @[LoadQueue.scala 141:18:@11938.4]
  wire  entriesToCheck_8_14; // @[LoadQueue.scala 141:26:@11939.4]
  wire  _T_13096; // @[LoadQueue.scala 141:18:@11940.4]
  wire  entriesToCheck_8_15; // @[LoadQueue.scala 141:26:@11941.4]
  wire  _T_13098; // @[LoadQueue.scala 141:18:@11958.4]
  wire  entriesToCheck_9_0; // @[LoadQueue.scala 141:26:@11959.4]
  wire  _T_13100; // @[LoadQueue.scala 141:18:@11960.4]
  wire  entriesToCheck_9_1; // @[LoadQueue.scala 141:26:@11961.4]
  wire  _T_13102; // @[LoadQueue.scala 141:18:@11962.4]
  wire  entriesToCheck_9_2; // @[LoadQueue.scala 141:26:@11963.4]
  wire  _T_13104; // @[LoadQueue.scala 141:18:@11964.4]
  wire  entriesToCheck_9_3; // @[LoadQueue.scala 141:26:@11965.4]
  wire  _T_13106; // @[LoadQueue.scala 141:18:@11966.4]
  wire  entriesToCheck_9_4; // @[LoadQueue.scala 141:26:@11967.4]
  wire  _T_13108; // @[LoadQueue.scala 141:18:@11968.4]
  wire  entriesToCheck_9_5; // @[LoadQueue.scala 141:26:@11969.4]
  wire  _T_13110; // @[LoadQueue.scala 141:18:@11970.4]
  wire  entriesToCheck_9_6; // @[LoadQueue.scala 141:26:@11971.4]
  wire  _T_13112; // @[LoadQueue.scala 141:18:@11972.4]
  wire  entriesToCheck_9_7; // @[LoadQueue.scala 141:26:@11973.4]
  wire  _T_13114; // @[LoadQueue.scala 141:18:@11974.4]
  wire  entriesToCheck_9_8; // @[LoadQueue.scala 141:26:@11975.4]
  wire  _T_13116; // @[LoadQueue.scala 141:18:@11976.4]
  wire  entriesToCheck_9_9; // @[LoadQueue.scala 141:26:@11977.4]
  wire  _T_13118; // @[LoadQueue.scala 141:18:@11978.4]
  wire  entriesToCheck_9_10; // @[LoadQueue.scala 141:26:@11979.4]
  wire  _T_13120; // @[LoadQueue.scala 141:18:@11980.4]
  wire  entriesToCheck_9_11; // @[LoadQueue.scala 141:26:@11981.4]
  wire  _T_13122; // @[LoadQueue.scala 141:18:@11982.4]
  wire  entriesToCheck_9_12; // @[LoadQueue.scala 141:26:@11983.4]
  wire  _T_13124; // @[LoadQueue.scala 141:18:@11984.4]
  wire  entriesToCheck_9_13; // @[LoadQueue.scala 141:26:@11985.4]
  wire  _T_13126; // @[LoadQueue.scala 141:18:@11986.4]
  wire  entriesToCheck_9_14; // @[LoadQueue.scala 141:26:@11987.4]
  wire  _T_13128; // @[LoadQueue.scala 141:18:@11988.4]
  wire  entriesToCheck_9_15; // @[LoadQueue.scala 141:26:@11989.4]
  wire  _T_13130; // @[LoadQueue.scala 141:18:@12006.4]
  wire  entriesToCheck_10_0; // @[LoadQueue.scala 141:26:@12007.4]
  wire  _T_13132; // @[LoadQueue.scala 141:18:@12008.4]
  wire  entriesToCheck_10_1; // @[LoadQueue.scala 141:26:@12009.4]
  wire  _T_13134; // @[LoadQueue.scala 141:18:@12010.4]
  wire  entriesToCheck_10_2; // @[LoadQueue.scala 141:26:@12011.4]
  wire  _T_13136; // @[LoadQueue.scala 141:18:@12012.4]
  wire  entriesToCheck_10_3; // @[LoadQueue.scala 141:26:@12013.4]
  wire  _T_13138; // @[LoadQueue.scala 141:18:@12014.4]
  wire  entriesToCheck_10_4; // @[LoadQueue.scala 141:26:@12015.4]
  wire  _T_13140; // @[LoadQueue.scala 141:18:@12016.4]
  wire  entriesToCheck_10_5; // @[LoadQueue.scala 141:26:@12017.4]
  wire  _T_13142; // @[LoadQueue.scala 141:18:@12018.4]
  wire  entriesToCheck_10_6; // @[LoadQueue.scala 141:26:@12019.4]
  wire  _T_13144; // @[LoadQueue.scala 141:18:@12020.4]
  wire  entriesToCheck_10_7; // @[LoadQueue.scala 141:26:@12021.4]
  wire  _T_13146; // @[LoadQueue.scala 141:18:@12022.4]
  wire  entriesToCheck_10_8; // @[LoadQueue.scala 141:26:@12023.4]
  wire  _T_13148; // @[LoadQueue.scala 141:18:@12024.4]
  wire  entriesToCheck_10_9; // @[LoadQueue.scala 141:26:@12025.4]
  wire  _T_13150; // @[LoadQueue.scala 141:18:@12026.4]
  wire  entriesToCheck_10_10; // @[LoadQueue.scala 141:26:@12027.4]
  wire  _T_13152; // @[LoadQueue.scala 141:18:@12028.4]
  wire  entriesToCheck_10_11; // @[LoadQueue.scala 141:26:@12029.4]
  wire  _T_13154; // @[LoadQueue.scala 141:18:@12030.4]
  wire  entriesToCheck_10_12; // @[LoadQueue.scala 141:26:@12031.4]
  wire  _T_13156; // @[LoadQueue.scala 141:18:@12032.4]
  wire  entriesToCheck_10_13; // @[LoadQueue.scala 141:26:@12033.4]
  wire  _T_13158; // @[LoadQueue.scala 141:18:@12034.4]
  wire  entriesToCheck_10_14; // @[LoadQueue.scala 141:26:@12035.4]
  wire  _T_13160; // @[LoadQueue.scala 141:18:@12036.4]
  wire  entriesToCheck_10_15; // @[LoadQueue.scala 141:26:@12037.4]
  wire  _T_13162; // @[LoadQueue.scala 141:18:@12054.4]
  wire  entriesToCheck_11_0; // @[LoadQueue.scala 141:26:@12055.4]
  wire  _T_13164; // @[LoadQueue.scala 141:18:@12056.4]
  wire  entriesToCheck_11_1; // @[LoadQueue.scala 141:26:@12057.4]
  wire  _T_13166; // @[LoadQueue.scala 141:18:@12058.4]
  wire  entriesToCheck_11_2; // @[LoadQueue.scala 141:26:@12059.4]
  wire  _T_13168; // @[LoadQueue.scala 141:18:@12060.4]
  wire  entriesToCheck_11_3; // @[LoadQueue.scala 141:26:@12061.4]
  wire  _T_13170; // @[LoadQueue.scala 141:18:@12062.4]
  wire  entriesToCheck_11_4; // @[LoadQueue.scala 141:26:@12063.4]
  wire  _T_13172; // @[LoadQueue.scala 141:18:@12064.4]
  wire  entriesToCheck_11_5; // @[LoadQueue.scala 141:26:@12065.4]
  wire  _T_13174; // @[LoadQueue.scala 141:18:@12066.4]
  wire  entriesToCheck_11_6; // @[LoadQueue.scala 141:26:@12067.4]
  wire  _T_13176; // @[LoadQueue.scala 141:18:@12068.4]
  wire  entriesToCheck_11_7; // @[LoadQueue.scala 141:26:@12069.4]
  wire  _T_13178; // @[LoadQueue.scala 141:18:@12070.4]
  wire  entriesToCheck_11_8; // @[LoadQueue.scala 141:26:@12071.4]
  wire  _T_13180; // @[LoadQueue.scala 141:18:@12072.4]
  wire  entriesToCheck_11_9; // @[LoadQueue.scala 141:26:@12073.4]
  wire  _T_13182; // @[LoadQueue.scala 141:18:@12074.4]
  wire  entriesToCheck_11_10; // @[LoadQueue.scala 141:26:@12075.4]
  wire  _T_13184; // @[LoadQueue.scala 141:18:@12076.4]
  wire  entriesToCheck_11_11; // @[LoadQueue.scala 141:26:@12077.4]
  wire  _T_13186; // @[LoadQueue.scala 141:18:@12078.4]
  wire  entriesToCheck_11_12; // @[LoadQueue.scala 141:26:@12079.4]
  wire  _T_13188; // @[LoadQueue.scala 141:18:@12080.4]
  wire  entriesToCheck_11_13; // @[LoadQueue.scala 141:26:@12081.4]
  wire  _T_13190; // @[LoadQueue.scala 141:18:@12082.4]
  wire  entriesToCheck_11_14; // @[LoadQueue.scala 141:26:@12083.4]
  wire  _T_13192; // @[LoadQueue.scala 141:18:@12084.4]
  wire  entriesToCheck_11_15; // @[LoadQueue.scala 141:26:@12085.4]
  wire  _T_13194; // @[LoadQueue.scala 141:18:@12102.4]
  wire  entriesToCheck_12_0; // @[LoadQueue.scala 141:26:@12103.4]
  wire  _T_13196; // @[LoadQueue.scala 141:18:@12104.4]
  wire  entriesToCheck_12_1; // @[LoadQueue.scala 141:26:@12105.4]
  wire  _T_13198; // @[LoadQueue.scala 141:18:@12106.4]
  wire  entriesToCheck_12_2; // @[LoadQueue.scala 141:26:@12107.4]
  wire  _T_13200; // @[LoadQueue.scala 141:18:@12108.4]
  wire  entriesToCheck_12_3; // @[LoadQueue.scala 141:26:@12109.4]
  wire  _T_13202; // @[LoadQueue.scala 141:18:@12110.4]
  wire  entriesToCheck_12_4; // @[LoadQueue.scala 141:26:@12111.4]
  wire  _T_13204; // @[LoadQueue.scala 141:18:@12112.4]
  wire  entriesToCheck_12_5; // @[LoadQueue.scala 141:26:@12113.4]
  wire  _T_13206; // @[LoadQueue.scala 141:18:@12114.4]
  wire  entriesToCheck_12_6; // @[LoadQueue.scala 141:26:@12115.4]
  wire  _T_13208; // @[LoadQueue.scala 141:18:@12116.4]
  wire  entriesToCheck_12_7; // @[LoadQueue.scala 141:26:@12117.4]
  wire  _T_13210; // @[LoadQueue.scala 141:18:@12118.4]
  wire  entriesToCheck_12_8; // @[LoadQueue.scala 141:26:@12119.4]
  wire  _T_13212; // @[LoadQueue.scala 141:18:@12120.4]
  wire  entriesToCheck_12_9; // @[LoadQueue.scala 141:26:@12121.4]
  wire  _T_13214; // @[LoadQueue.scala 141:18:@12122.4]
  wire  entriesToCheck_12_10; // @[LoadQueue.scala 141:26:@12123.4]
  wire  _T_13216; // @[LoadQueue.scala 141:18:@12124.4]
  wire  entriesToCheck_12_11; // @[LoadQueue.scala 141:26:@12125.4]
  wire  _T_13218; // @[LoadQueue.scala 141:18:@12126.4]
  wire  entriesToCheck_12_12; // @[LoadQueue.scala 141:26:@12127.4]
  wire  _T_13220; // @[LoadQueue.scala 141:18:@12128.4]
  wire  entriesToCheck_12_13; // @[LoadQueue.scala 141:26:@12129.4]
  wire  _T_13222; // @[LoadQueue.scala 141:18:@12130.4]
  wire  entriesToCheck_12_14; // @[LoadQueue.scala 141:26:@12131.4]
  wire  _T_13224; // @[LoadQueue.scala 141:18:@12132.4]
  wire  entriesToCheck_12_15; // @[LoadQueue.scala 141:26:@12133.4]
  wire  _T_13226; // @[LoadQueue.scala 141:18:@12150.4]
  wire  entriesToCheck_13_0; // @[LoadQueue.scala 141:26:@12151.4]
  wire  _T_13228; // @[LoadQueue.scala 141:18:@12152.4]
  wire  entriesToCheck_13_1; // @[LoadQueue.scala 141:26:@12153.4]
  wire  _T_13230; // @[LoadQueue.scala 141:18:@12154.4]
  wire  entriesToCheck_13_2; // @[LoadQueue.scala 141:26:@12155.4]
  wire  _T_13232; // @[LoadQueue.scala 141:18:@12156.4]
  wire  entriesToCheck_13_3; // @[LoadQueue.scala 141:26:@12157.4]
  wire  _T_13234; // @[LoadQueue.scala 141:18:@12158.4]
  wire  entriesToCheck_13_4; // @[LoadQueue.scala 141:26:@12159.4]
  wire  _T_13236; // @[LoadQueue.scala 141:18:@12160.4]
  wire  entriesToCheck_13_5; // @[LoadQueue.scala 141:26:@12161.4]
  wire  _T_13238; // @[LoadQueue.scala 141:18:@12162.4]
  wire  entriesToCheck_13_6; // @[LoadQueue.scala 141:26:@12163.4]
  wire  _T_13240; // @[LoadQueue.scala 141:18:@12164.4]
  wire  entriesToCheck_13_7; // @[LoadQueue.scala 141:26:@12165.4]
  wire  _T_13242; // @[LoadQueue.scala 141:18:@12166.4]
  wire  entriesToCheck_13_8; // @[LoadQueue.scala 141:26:@12167.4]
  wire  _T_13244; // @[LoadQueue.scala 141:18:@12168.4]
  wire  entriesToCheck_13_9; // @[LoadQueue.scala 141:26:@12169.4]
  wire  _T_13246; // @[LoadQueue.scala 141:18:@12170.4]
  wire  entriesToCheck_13_10; // @[LoadQueue.scala 141:26:@12171.4]
  wire  _T_13248; // @[LoadQueue.scala 141:18:@12172.4]
  wire  entriesToCheck_13_11; // @[LoadQueue.scala 141:26:@12173.4]
  wire  _T_13250; // @[LoadQueue.scala 141:18:@12174.4]
  wire  entriesToCheck_13_12; // @[LoadQueue.scala 141:26:@12175.4]
  wire  _T_13252; // @[LoadQueue.scala 141:18:@12176.4]
  wire  entriesToCheck_13_13; // @[LoadQueue.scala 141:26:@12177.4]
  wire  _T_13254; // @[LoadQueue.scala 141:18:@12178.4]
  wire  entriesToCheck_13_14; // @[LoadQueue.scala 141:26:@12179.4]
  wire  _T_13256; // @[LoadQueue.scala 141:18:@12180.4]
  wire  entriesToCheck_13_15; // @[LoadQueue.scala 141:26:@12181.4]
  wire  _T_13258; // @[LoadQueue.scala 141:18:@12198.4]
  wire  entriesToCheck_14_0; // @[LoadQueue.scala 141:26:@12199.4]
  wire  _T_13260; // @[LoadQueue.scala 141:18:@12200.4]
  wire  entriesToCheck_14_1; // @[LoadQueue.scala 141:26:@12201.4]
  wire  _T_13262; // @[LoadQueue.scala 141:18:@12202.4]
  wire  entriesToCheck_14_2; // @[LoadQueue.scala 141:26:@12203.4]
  wire  _T_13264; // @[LoadQueue.scala 141:18:@12204.4]
  wire  entriesToCheck_14_3; // @[LoadQueue.scala 141:26:@12205.4]
  wire  _T_13266; // @[LoadQueue.scala 141:18:@12206.4]
  wire  entriesToCheck_14_4; // @[LoadQueue.scala 141:26:@12207.4]
  wire  _T_13268; // @[LoadQueue.scala 141:18:@12208.4]
  wire  entriesToCheck_14_5; // @[LoadQueue.scala 141:26:@12209.4]
  wire  _T_13270; // @[LoadQueue.scala 141:18:@12210.4]
  wire  entriesToCheck_14_6; // @[LoadQueue.scala 141:26:@12211.4]
  wire  _T_13272; // @[LoadQueue.scala 141:18:@12212.4]
  wire  entriesToCheck_14_7; // @[LoadQueue.scala 141:26:@12213.4]
  wire  _T_13274; // @[LoadQueue.scala 141:18:@12214.4]
  wire  entriesToCheck_14_8; // @[LoadQueue.scala 141:26:@12215.4]
  wire  _T_13276; // @[LoadQueue.scala 141:18:@12216.4]
  wire  entriesToCheck_14_9; // @[LoadQueue.scala 141:26:@12217.4]
  wire  _T_13278; // @[LoadQueue.scala 141:18:@12218.4]
  wire  entriesToCheck_14_10; // @[LoadQueue.scala 141:26:@12219.4]
  wire  _T_13280; // @[LoadQueue.scala 141:18:@12220.4]
  wire  entriesToCheck_14_11; // @[LoadQueue.scala 141:26:@12221.4]
  wire  _T_13282; // @[LoadQueue.scala 141:18:@12222.4]
  wire  entriesToCheck_14_12; // @[LoadQueue.scala 141:26:@12223.4]
  wire  _T_13284; // @[LoadQueue.scala 141:18:@12224.4]
  wire  entriesToCheck_14_13; // @[LoadQueue.scala 141:26:@12225.4]
  wire  _T_13286; // @[LoadQueue.scala 141:18:@12226.4]
  wire  entriesToCheck_14_14; // @[LoadQueue.scala 141:26:@12227.4]
  wire  _T_13288; // @[LoadQueue.scala 141:18:@12228.4]
  wire  entriesToCheck_14_15; // @[LoadQueue.scala 141:26:@12229.4]
  wire  _T_13290; // @[LoadQueue.scala 141:18:@12246.4]
  wire  entriesToCheck_15_0; // @[LoadQueue.scala 141:26:@12247.4]
  wire  _T_13292; // @[LoadQueue.scala 141:18:@12248.4]
  wire  entriesToCheck_15_1; // @[LoadQueue.scala 141:26:@12249.4]
  wire  _T_13294; // @[LoadQueue.scala 141:18:@12250.4]
  wire  entriesToCheck_15_2; // @[LoadQueue.scala 141:26:@12251.4]
  wire  _T_13296; // @[LoadQueue.scala 141:18:@12252.4]
  wire  entriesToCheck_15_3; // @[LoadQueue.scala 141:26:@12253.4]
  wire  _T_13298; // @[LoadQueue.scala 141:18:@12254.4]
  wire  entriesToCheck_15_4; // @[LoadQueue.scala 141:26:@12255.4]
  wire  _T_13300; // @[LoadQueue.scala 141:18:@12256.4]
  wire  entriesToCheck_15_5; // @[LoadQueue.scala 141:26:@12257.4]
  wire  _T_13302; // @[LoadQueue.scala 141:18:@12258.4]
  wire  entriesToCheck_15_6; // @[LoadQueue.scala 141:26:@12259.4]
  wire  _T_13304; // @[LoadQueue.scala 141:18:@12260.4]
  wire  entriesToCheck_15_7; // @[LoadQueue.scala 141:26:@12261.4]
  wire  _T_13306; // @[LoadQueue.scala 141:18:@12262.4]
  wire  entriesToCheck_15_8; // @[LoadQueue.scala 141:26:@12263.4]
  wire  _T_13308; // @[LoadQueue.scala 141:18:@12264.4]
  wire  entriesToCheck_15_9; // @[LoadQueue.scala 141:26:@12265.4]
  wire  _T_13310; // @[LoadQueue.scala 141:18:@12266.4]
  wire  entriesToCheck_15_10; // @[LoadQueue.scala 141:26:@12267.4]
  wire  _T_13312; // @[LoadQueue.scala 141:18:@12268.4]
  wire  entriesToCheck_15_11; // @[LoadQueue.scala 141:26:@12269.4]
  wire  _T_13314; // @[LoadQueue.scala 141:18:@12270.4]
  wire  entriesToCheck_15_12; // @[LoadQueue.scala 141:26:@12271.4]
  wire  _T_13316; // @[LoadQueue.scala 141:18:@12272.4]
  wire  entriesToCheck_15_13; // @[LoadQueue.scala 141:26:@12273.4]
  wire  _T_13318; // @[LoadQueue.scala 141:18:@12274.4]
  wire  entriesToCheck_15_14; // @[LoadQueue.scala 141:26:@12275.4]
  wire  _T_13320; // @[LoadQueue.scala 141:18:@12276.4]
  wire  entriesToCheck_15_15; // @[LoadQueue.scala 141:26:@12277.4]
  wire  _T_14552; // @[LoadQueue.scala 151:92:@12295.4]
  wire  _T_14553; // @[LoadQueue.scala 152:41:@12296.4]
  wire  _T_14554; // @[LoadQueue.scala 153:30:@12297.4]
  wire  conflict_0_0; // @[LoadQueue.scala 152:68:@12298.4]
  wire  _T_14556; // @[LoadQueue.scala 151:92:@12300.4]
  wire  _T_14557; // @[LoadQueue.scala 152:41:@12301.4]
  wire  _T_14558; // @[LoadQueue.scala 153:30:@12302.4]
  wire  conflict_0_1; // @[LoadQueue.scala 152:68:@12303.4]
  wire  _T_14560; // @[LoadQueue.scala 151:92:@12305.4]
  wire  _T_14561; // @[LoadQueue.scala 152:41:@12306.4]
  wire  _T_14562; // @[LoadQueue.scala 153:30:@12307.4]
  wire  conflict_0_2; // @[LoadQueue.scala 152:68:@12308.4]
  wire  _T_14564; // @[LoadQueue.scala 151:92:@12310.4]
  wire  _T_14565; // @[LoadQueue.scala 152:41:@12311.4]
  wire  _T_14566; // @[LoadQueue.scala 153:30:@12312.4]
  wire  conflict_0_3; // @[LoadQueue.scala 152:68:@12313.4]
  wire  _T_14568; // @[LoadQueue.scala 151:92:@12315.4]
  wire  _T_14569; // @[LoadQueue.scala 152:41:@12316.4]
  wire  _T_14570; // @[LoadQueue.scala 153:30:@12317.4]
  wire  conflict_0_4; // @[LoadQueue.scala 152:68:@12318.4]
  wire  _T_14572; // @[LoadQueue.scala 151:92:@12320.4]
  wire  _T_14573; // @[LoadQueue.scala 152:41:@12321.4]
  wire  _T_14574; // @[LoadQueue.scala 153:30:@12322.4]
  wire  conflict_0_5; // @[LoadQueue.scala 152:68:@12323.4]
  wire  _T_14576; // @[LoadQueue.scala 151:92:@12325.4]
  wire  _T_14577; // @[LoadQueue.scala 152:41:@12326.4]
  wire  _T_14578; // @[LoadQueue.scala 153:30:@12327.4]
  wire  conflict_0_6; // @[LoadQueue.scala 152:68:@12328.4]
  wire  _T_14580; // @[LoadQueue.scala 151:92:@12330.4]
  wire  _T_14581; // @[LoadQueue.scala 152:41:@12331.4]
  wire  _T_14582; // @[LoadQueue.scala 153:30:@12332.4]
  wire  conflict_0_7; // @[LoadQueue.scala 152:68:@12333.4]
  wire  _T_14584; // @[LoadQueue.scala 151:92:@12335.4]
  wire  _T_14585; // @[LoadQueue.scala 152:41:@12336.4]
  wire  _T_14586; // @[LoadQueue.scala 153:30:@12337.4]
  wire  conflict_0_8; // @[LoadQueue.scala 152:68:@12338.4]
  wire  _T_14588; // @[LoadQueue.scala 151:92:@12340.4]
  wire  _T_14589; // @[LoadQueue.scala 152:41:@12341.4]
  wire  _T_14590; // @[LoadQueue.scala 153:30:@12342.4]
  wire  conflict_0_9; // @[LoadQueue.scala 152:68:@12343.4]
  wire  _T_14592; // @[LoadQueue.scala 151:92:@12345.4]
  wire  _T_14593; // @[LoadQueue.scala 152:41:@12346.4]
  wire  _T_14594; // @[LoadQueue.scala 153:30:@12347.4]
  wire  conflict_0_10; // @[LoadQueue.scala 152:68:@12348.4]
  wire  _T_14596; // @[LoadQueue.scala 151:92:@12350.4]
  wire  _T_14597; // @[LoadQueue.scala 152:41:@12351.4]
  wire  _T_14598; // @[LoadQueue.scala 153:30:@12352.4]
  wire  conflict_0_11; // @[LoadQueue.scala 152:68:@12353.4]
  wire  _T_14600; // @[LoadQueue.scala 151:92:@12355.4]
  wire  _T_14601; // @[LoadQueue.scala 152:41:@12356.4]
  wire  _T_14602; // @[LoadQueue.scala 153:30:@12357.4]
  wire  conflict_0_12; // @[LoadQueue.scala 152:68:@12358.4]
  wire  _T_14604; // @[LoadQueue.scala 151:92:@12360.4]
  wire  _T_14605; // @[LoadQueue.scala 152:41:@12361.4]
  wire  _T_14606; // @[LoadQueue.scala 153:30:@12362.4]
  wire  conflict_0_13; // @[LoadQueue.scala 152:68:@12363.4]
  wire  _T_14608; // @[LoadQueue.scala 151:92:@12365.4]
  wire  _T_14609; // @[LoadQueue.scala 152:41:@12366.4]
  wire  _T_14610; // @[LoadQueue.scala 153:30:@12367.4]
  wire  conflict_0_14; // @[LoadQueue.scala 152:68:@12368.4]
  wire  _T_14612; // @[LoadQueue.scala 151:92:@12370.4]
  wire  _T_14613; // @[LoadQueue.scala 152:41:@12371.4]
  wire  _T_14614; // @[LoadQueue.scala 153:30:@12372.4]
  wire  conflict_0_15; // @[LoadQueue.scala 152:68:@12373.4]
  wire  _T_14616; // @[LoadQueue.scala 151:92:@12375.4]
  wire  _T_14617; // @[LoadQueue.scala 152:41:@12376.4]
  wire  _T_14618; // @[LoadQueue.scala 153:30:@12377.4]
  wire  conflict_1_0; // @[LoadQueue.scala 152:68:@12378.4]
  wire  _T_14620; // @[LoadQueue.scala 151:92:@12380.4]
  wire  _T_14621; // @[LoadQueue.scala 152:41:@12381.4]
  wire  _T_14622; // @[LoadQueue.scala 153:30:@12382.4]
  wire  conflict_1_1; // @[LoadQueue.scala 152:68:@12383.4]
  wire  _T_14624; // @[LoadQueue.scala 151:92:@12385.4]
  wire  _T_14625; // @[LoadQueue.scala 152:41:@12386.4]
  wire  _T_14626; // @[LoadQueue.scala 153:30:@12387.4]
  wire  conflict_1_2; // @[LoadQueue.scala 152:68:@12388.4]
  wire  _T_14628; // @[LoadQueue.scala 151:92:@12390.4]
  wire  _T_14629; // @[LoadQueue.scala 152:41:@12391.4]
  wire  _T_14630; // @[LoadQueue.scala 153:30:@12392.4]
  wire  conflict_1_3; // @[LoadQueue.scala 152:68:@12393.4]
  wire  _T_14632; // @[LoadQueue.scala 151:92:@12395.4]
  wire  _T_14633; // @[LoadQueue.scala 152:41:@12396.4]
  wire  _T_14634; // @[LoadQueue.scala 153:30:@12397.4]
  wire  conflict_1_4; // @[LoadQueue.scala 152:68:@12398.4]
  wire  _T_14636; // @[LoadQueue.scala 151:92:@12400.4]
  wire  _T_14637; // @[LoadQueue.scala 152:41:@12401.4]
  wire  _T_14638; // @[LoadQueue.scala 153:30:@12402.4]
  wire  conflict_1_5; // @[LoadQueue.scala 152:68:@12403.4]
  wire  _T_14640; // @[LoadQueue.scala 151:92:@12405.4]
  wire  _T_14641; // @[LoadQueue.scala 152:41:@12406.4]
  wire  _T_14642; // @[LoadQueue.scala 153:30:@12407.4]
  wire  conflict_1_6; // @[LoadQueue.scala 152:68:@12408.4]
  wire  _T_14644; // @[LoadQueue.scala 151:92:@12410.4]
  wire  _T_14645; // @[LoadQueue.scala 152:41:@12411.4]
  wire  _T_14646; // @[LoadQueue.scala 153:30:@12412.4]
  wire  conflict_1_7; // @[LoadQueue.scala 152:68:@12413.4]
  wire  _T_14648; // @[LoadQueue.scala 151:92:@12415.4]
  wire  _T_14649; // @[LoadQueue.scala 152:41:@12416.4]
  wire  _T_14650; // @[LoadQueue.scala 153:30:@12417.4]
  wire  conflict_1_8; // @[LoadQueue.scala 152:68:@12418.4]
  wire  _T_14652; // @[LoadQueue.scala 151:92:@12420.4]
  wire  _T_14653; // @[LoadQueue.scala 152:41:@12421.4]
  wire  _T_14654; // @[LoadQueue.scala 153:30:@12422.4]
  wire  conflict_1_9; // @[LoadQueue.scala 152:68:@12423.4]
  wire  _T_14656; // @[LoadQueue.scala 151:92:@12425.4]
  wire  _T_14657; // @[LoadQueue.scala 152:41:@12426.4]
  wire  _T_14658; // @[LoadQueue.scala 153:30:@12427.4]
  wire  conflict_1_10; // @[LoadQueue.scala 152:68:@12428.4]
  wire  _T_14660; // @[LoadQueue.scala 151:92:@12430.4]
  wire  _T_14661; // @[LoadQueue.scala 152:41:@12431.4]
  wire  _T_14662; // @[LoadQueue.scala 153:30:@12432.4]
  wire  conflict_1_11; // @[LoadQueue.scala 152:68:@12433.4]
  wire  _T_14664; // @[LoadQueue.scala 151:92:@12435.4]
  wire  _T_14665; // @[LoadQueue.scala 152:41:@12436.4]
  wire  _T_14666; // @[LoadQueue.scala 153:30:@12437.4]
  wire  conflict_1_12; // @[LoadQueue.scala 152:68:@12438.4]
  wire  _T_14668; // @[LoadQueue.scala 151:92:@12440.4]
  wire  _T_14669; // @[LoadQueue.scala 152:41:@12441.4]
  wire  _T_14670; // @[LoadQueue.scala 153:30:@12442.4]
  wire  conflict_1_13; // @[LoadQueue.scala 152:68:@12443.4]
  wire  _T_14672; // @[LoadQueue.scala 151:92:@12445.4]
  wire  _T_14673; // @[LoadQueue.scala 152:41:@12446.4]
  wire  _T_14674; // @[LoadQueue.scala 153:30:@12447.4]
  wire  conflict_1_14; // @[LoadQueue.scala 152:68:@12448.4]
  wire  _T_14676; // @[LoadQueue.scala 151:92:@12450.4]
  wire  _T_14677; // @[LoadQueue.scala 152:41:@12451.4]
  wire  _T_14678; // @[LoadQueue.scala 153:30:@12452.4]
  wire  conflict_1_15; // @[LoadQueue.scala 152:68:@12453.4]
  wire  _T_14680; // @[LoadQueue.scala 151:92:@12455.4]
  wire  _T_14681; // @[LoadQueue.scala 152:41:@12456.4]
  wire  _T_14682; // @[LoadQueue.scala 153:30:@12457.4]
  wire  conflict_2_0; // @[LoadQueue.scala 152:68:@12458.4]
  wire  _T_14684; // @[LoadQueue.scala 151:92:@12460.4]
  wire  _T_14685; // @[LoadQueue.scala 152:41:@12461.4]
  wire  _T_14686; // @[LoadQueue.scala 153:30:@12462.4]
  wire  conflict_2_1; // @[LoadQueue.scala 152:68:@12463.4]
  wire  _T_14688; // @[LoadQueue.scala 151:92:@12465.4]
  wire  _T_14689; // @[LoadQueue.scala 152:41:@12466.4]
  wire  _T_14690; // @[LoadQueue.scala 153:30:@12467.4]
  wire  conflict_2_2; // @[LoadQueue.scala 152:68:@12468.4]
  wire  _T_14692; // @[LoadQueue.scala 151:92:@12470.4]
  wire  _T_14693; // @[LoadQueue.scala 152:41:@12471.4]
  wire  _T_14694; // @[LoadQueue.scala 153:30:@12472.4]
  wire  conflict_2_3; // @[LoadQueue.scala 152:68:@12473.4]
  wire  _T_14696; // @[LoadQueue.scala 151:92:@12475.4]
  wire  _T_14697; // @[LoadQueue.scala 152:41:@12476.4]
  wire  _T_14698; // @[LoadQueue.scala 153:30:@12477.4]
  wire  conflict_2_4; // @[LoadQueue.scala 152:68:@12478.4]
  wire  _T_14700; // @[LoadQueue.scala 151:92:@12480.4]
  wire  _T_14701; // @[LoadQueue.scala 152:41:@12481.4]
  wire  _T_14702; // @[LoadQueue.scala 153:30:@12482.4]
  wire  conflict_2_5; // @[LoadQueue.scala 152:68:@12483.4]
  wire  _T_14704; // @[LoadQueue.scala 151:92:@12485.4]
  wire  _T_14705; // @[LoadQueue.scala 152:41:@12486.4]
  wire  _T_14706; // @[LoadQueue.scala 153:30:@12487.4]
  wire  conflict_2_6; // @[LoadQueue.scala 152:68:@12488.4]
  wire  _T_14708; // @[LoadQueue.scala 151:92:@12490.4]
  wire  _T_14709; // @[LoadQueue.scala 152:41:@12491.4]
  wire  _T_14710; // @[LoadQueue.scala 153:30:@12492.4]
  wire  conflict_2_7; // @[LoadQueue.scala 152:68:@12493.4]
  wire  _T_14712; // @[LoadQueue.scala 151:92:@12495.4]
  wire  _T_14713; // @[LoadQueue.scala 152:41:@12496.4]
  wire  _T_14714; // @[LoadQueue.scala 153:30:@12497.4]
  wire  conflict_2_8; // @[LoadQueue.scala 152:68:@12498.4]
  wire  _T_14716; // @[LoadQueue.scala 151:92:@12500.4]
  wire  _T_14717; // @[LoadQueue.scala 152:41:@12501.4]
  wire  _T_14718; // @[LoadQueue.scala 153:30:@12502.4]
  wire  conflict_2_9; // @[LoadQueue.scala 152:68:@12503.4]
  wire  _T_14720; // @[LoadQueue.scala 151:92:@12505.4]
  wire  _T_14721; // @[LoadQueue.scala 152:41:@12506.4]
  wire  _T_14722; // @[LoadQueue.scala 153:30:@12507.4]
  wire  conflict_2_10; // @[LoadQueue.scala 152:68:@12508.4]
  wire  _T_14724; // @[LoadQueue.scala 151:92:@12510.4]
  wire  _T_14725; // @[LoadQueue.scala 152:41:@12511.4]
  wire  _T_14726; // @[LoadQueue.scala 153:30:@12512.4]
  wire  conflict_2_11; // @[LoadQueue.scala 152:68:@12513.4]
  wire  _T_14728; // @[LoadQueue.scala 151:92:@12515.4]
  wire  _T_14729; // @[LoadQueue.scala 152:41:@12516.4]
  wire  _T_14730; // @[LoadQueue.scala 153:30:@12517.4]
  wire  conflict_2_12; // @[LoadQueue.scala 152:68:@12518.4]
  wire  _T_14732; // @[LoadQueue.scala 151:92:@12520.4]
  wire  _T_14733; // @[LoadQueue.scala 152:41:@12521.4]
  wire  _T_14734; // @[LoadQueue.scala 153:30:@12522.4]
  wire  conflict_2_13; // @[LoadQueue.scala 152:68:@12523.4]
  wire  _T_14736; // @[LoadQueue.scala 151:92:@12525.4]
  wire  _T_14737; // @[LoadQueue.scala 152:41:@12526.4]
  wire  _T_14738; // @[LoadQueue.scala 153:30:@12527.4]
  wire  conflict_2_14; // @[LoadQueue.scala 152:68:@12528.4]
  wire  _T_14740; // @[LoadQueue.scala 151:92:@12530.4]
  wire  _T_14741; // @[LoadQueue.scala 152:41:@12531.4]
  wire  _T_14742; // @[LoadQueue.scala 153:30:@12532.4]
  wire  conflict_2_15; // @[LoadQueue.scala 152:68:@12533.4]
  wire  _T_14744; // @[LoadQueue.scala 151:92:@12535.4]
  wire  _T_14745; // @[LoadQueue.scala 152:41:@12536.4]
  wire  _T_14746; // @[LoadQueue.scala 153:30:@12537.4]
  wire  conflict_3_0; // @[LoadQueue.scala 152:68:@12538.4]
  wire  _T_14748; // @[LoadQueue.scala 151:92:@12540.4]
  wire  _T_14749; // @[LoadQueue.scala 152:41:@12541.4]
  wire  _T_14750; // @[LoadQueue.scala 153:30:@12542.4]
  wire  conflict_3_1; // @[LoadQueue.scala 152:68:@12543.4]
  wire  _T_14752; // @[LoadQueue.scala 151:92:@12545.4]
  wire  _T_14753; // @[LoadQueue.scala 152:41:@12546.4]
  wire  _T_14754; // @[LoadQueue.scala 153:30:@12547.4]
  wire  conflict_3_2; // @[LoadQueue.scala 152:68:@12548.4]
  wire  _T_14756; // @[LoadQueue.scala 151:92:@12550.4]
  wire  _T_14757; // @[LoadQueue.scala 152:41:@12551.4]
  wire  _T_14758; // @[LoadQueue.scala 153:30:@12552.4]
  wire  conflict_3_3; // @[LoadQueue.scala 152:68:@12553.4]
  wire  _T_14760; // @[LoadQueue.scala 151:92:@12555.4]
  wire  _T_14761; // @[LoadQueue.scala 152:41:@12556.4]
  wire  _T_14762; // @[LoadQueue.scala 153:30:@12557.4]
  wire  conflict_3_4; // @[LoadQueue.scala 152:68:@12558.4]
  wire  _T_14764; // @[LoadQueue.scala 151:92:@12560.4]
  wire  _T_14765; // @[LoadQueue.scala 152:41:@12561.4]
  wire  _T_14766; // @[LoadQueue.scala 153:30:@12562.4]
  wire  conflict_3_5; // @[LoadQueue.scala 152:68:@12563.4]
  wire  _T_14768; // @[LoadQueue.scala 151:92:@12565.4]
  wire  _T_14769; // @[LoadQueue.scala 152:41:@12566.4]
  wire  _T_14770; // @[LoadQueue.scala 153:30:@12567.4]
  wire  conflict_3_6; // @[LoadQueue.scala 152:68:@12568.4]
  wire  _T_14772; // @[LoadQueue.scala 151:92:@12570.4]
  wire  _T_14773; // @[LoadQueue.scala 152:41:@12571.4]
  wire  _T_14774; // @[LoadQueue.scala 153:30:@12572.4]
  wire  conflict_3_7; // @[LoadQueue.scala 152:68:@12573.4]
  wire  _T_14776; // @[LoadQueue.scala 151:92:@12575.4]
  wire  _T_14777; // @[LoadQueue.scala 152:41:@12576.4]
  wire  _T_14778; // @[LoadQueue.scala 153:30:@12577.4]
  wire  conflict_3_8; // @[LoadQueue.scala 152:68:@12578.4]
  wire  _T_14780; // @[LoadQueue.scala 151:92:@12580.4]
  wire  _T_14781; // @[LoadQueue.scala 152:41:@12581.4]
  wire  _T_14782; // @[LoadQueue.scala 153:30:@12582.4]
  wire  conflict_3_9; // @[LoadQueue.scala 152:68:@12583.4]
  wire  _T_14784; // @[LoadQueue.scala 151:92:@12585.4]
  wire  _T_14785; // @[LoadQueue.scala 152:41:@12586.4]
  wire  _T_14786; // @[LoadQueue.scala 153:30:@12587.4]
  wire  conflict_3_10; // @[LoadQueue.scala 152:68:@12588.4]
  wire  _T_14788; // @[LoadQueue.scala 151:92:@12590.4]
  wire  _T_14789; // @[LoadQueue.scala 152:41:@12591.4]
  wire  _T_14790; // @[LoadQueue.scala 153:30:@12592.4]
  wire  conflict_3_11; // @[LoadQueue.scala 152:68:@12593.4]
  wire  _T_14792; // @[LoadQueue.scala 151:92:@12595.4]
  wire  _T_14793; // @[LoadQueue.scala 152:41:@12596.4]
  wire  _T_14794; // @[LoadQueue.scala 153:30:@12597.4]
  wire  conflict_3_12; // @[LoadQueue.scala 152:68:@12598.4]
  wire  _T_14796; // @[LoadQueue.scala 151:92:@12600.4]
  wire  _T_14797; // @[LoadQueue.scala 152:41:@12601.4]
  wire  _T_14798; // @[LoadQueue.scala 153:30:@12602.4]
  wire  conflict_3_13; // @[LoadQueue.scala 152:68:@12603.4]
  wire  _T_14800; // @[LoadQueue.scala 151:92:@12605.4]
  wire  _T_14801; // @[LoadQueue.scala 152:41:@12606.4]
  wire  _T_14802; // @[LoadQueue.scala 153:30:@12607.4]
  wire  conflict_3_14; // @[LoadQueue.scala 152:68:@12608.4]
  wire  _T_14804; // @[LoadQueue.scala 151:92:@12610.4]
  wire  _T_14805; // @[LoadQueue.scala 152:41:@12611.4]
  wire  _T_14806; // @[LoadQueue.scala 153:30:@12612.4]
  wire  conflict_3_15; // @[LoadQueue.scala 152:68:@12613.4]
  wire  _T_14808; // @[LoadQueue.scala 151:92:@12615.4]
  wire  _T_14809; // @[LoadQueue.scala 152:41:@12616.4]
  wire  _T_14810; // @[LoadQueue.scala 153:30:@12617.4]
  wire  conflict_4_0; // @[LoadQueue.scala 152:68:@12618.4]
  wire  _T_14812; // @[LoadQueue.scala 151:92:@12620.4]
  wire  _T_14813; // @[LoadQueue.scala 152:41:@12621.4]
  wire  _T_14814; // @[LoadQueue.scala 153:30:@12622.4]
  wire  conflict_4_1; // @[LoadQueue.scala 152:68:@12623.4]
  wire  _T_14816; // @[LoadQueue.scala 151:92:@12625.4]
  wire  _T_14817; // @[LoadQueue.scala 152:41:@12626.4]
  wire  _T_14818; // @[LoadQueue.scala 153:30:@12627.4]
  wire  conflict_4_2; // @[LoadQueue.scala 152:68:@12628.4]
  wire  _T_14820; // @[LoadQueue.scala 151:92:@12630.4]
  wire  _T_14821; // @[LoadQueue.scala 152:41:@12631.4]
  wire  _T_14822; // @[LoadQueue.scala 153:30:@12632.4]
  wire  conflict_4_3; // @[LoadQueue.scala 152:68:@12633.4]
  wire  _T_14824; // @[LoadQueue.scala 151:92:@12635.4]
  wire  _T_14825; // @[LoadQueue.scala 152:41:@12636.4]
  wire  _T_14826; // @[LoadQueue.scala 153:30:@12637.4]
  wire  conflict_4_4; // @[LoadQueue.scala 152:68:@12638.4]
  wire  _T_14828; // @[LoadQueue.scala 151:92:@12640.4]
  wire  _T_14829; // @[LoadQueue.scala 152:41:@12641.4]
  wire  _T_14830; // @[LoadQueue.scala 153:30:@12642.4]
  wire  conflict_4_5; // @[LoadQueue.scala 152:68:@12643.4]
  wire  _T_14832; // @[LoadQueue.scala 151:92:@12645.4]
  wire  _T_14833; // @[LoadQueue.scala 152:41:@12646.4]
  wire  _T_14834; // @[LoadQueue.scala 153:30:@12647.4]
  wire  conflict_4_6; // @[LoadQueue.scala 152:68:@12648.4]
  wire  _T_14836; // @[LoadQueue.scala 151:92:@12650.4]
  wire  _T_14837; // @[LoadQueue.scala 152:41:@12651.4]
  wire  _T_14838; // @[LoadQueue.scala 153:30:@12652.4]
  wire  conflict_4_7; // @[LoadQueue.scala 152:68:@12653.4]
  wire  _T_14840; // @[LoadQueue.scala 151:92:@12655.4]
  wire  _T_14841; // @[LoadQueue.scala 152:41:@12656.4]
  wire  _T_14842; // @[LoadQueue.scala 153:30:@12657.4]
  wire  conflict_4_8; // @[LoadQueue.scala 152:68:@12658.4]
  wire  _T_14844; // @[LoadQueue.scala 151:92:@12660.4]
  wire  _T_14845; // @[LoadQueue.scala 152:41:@12661.4]
  wire  _T_14846; // @[LoadQueue.scala 153:30:@12662.4]
  wire  conflict_4_9; // @[LoadQueue.scala 152:68:@12663.4]
  wire  _T_14848; // @[LoadQueue.scala 151:92:@12665.4]
  wire  _T_14849; // @[LoadQueue.scala 152:41:@12666.4]
  wire  _T_14850; // @[LoadQueue.scala 153:30:@12667.4]
  wire  conflict_4_10; // @[LoadQueue.scala 152:68:@12668.4]
  wire  _T_14852; // @[LoadQueue.scala 151:92:@12670.4]
  wire  _T_14853; // @[LoadQueue.scala 152:41:@12671.4]
  wire  _T_14854; // @[LoadQueue.scala 153:30:@12672.4]
  wire  conflict_4_11; // @[LoadQueue.scala 152:68:@12673.4]
  wire  _T_14856; // @[LoadQueue.scala 151:92:@12675.4]
  wire  _T_14857; // @[LoadQueue.scala 152:41:@12676.4]
  wire  _T_14858; // @[LoadQueue.scala 153:30:@12677.4]
  wire  conflict_4_12; // @[LoadQueue.scala 152:68:@12678.4]
  wire  _T_14860; // @[LoadQueue.scala 151:92:@12680.4]
  wire  _T_14861; // @[LoadQueue.scala 152:41:@12681.4]
  wire  _T_14862; // @[LoadQueue.scala 153:30:@12682.4]
  wire  conflict_4_13; // @[LoadQueue.scala 152:68:@12683.4]
  wire  _T_14864; // @[LoadQueue.scala 151:92:@12685.4]
  wire  _T_14865; // @[LoadQueue.scala 152:41:@12686.4]
  wire  _T_14866; // @[LoadQueue.scala 153:30:@12687.4]
  wire  conflict_4_14; // @[LoadQueue.scala 152:68:@12688.4]
  wire  _T_14868; // @[LoadQueue.scala 151:92:@12690.4]
  wire  _T_14869; // @[LoadQueue.scala 152:41:@12691.4]
  wire  _T_14870; // @[LoadQueue.scala 153:30:@12692.4]
  wire  conflict_4_15; // @[LoadQueue.scala 152:68:@12693.4]
  wire  _T_14872; // @[LoadQueue.scala 151:92:@12695.4]
  wire  _T_14873; // @[LoadQueue.scala 152:41:@12696.4]
  wire  _T_14874; // @[LoadQueue.scala 153:30:@12697.4]
  wire  conflict_5_0; // @[LoadQueue.scala 152:68:@12698.4]
  wire  _T_14876; // @[LoadQueue.scala 151:92:@12700.4]
  wire  _T_14877; // @[LoadQueue.scala 152:41:@12701.4]
  wire  _T_14878; // @[LoadQueue.scala 153:30:@12702.4]
  wire  conflict_5_1; // @[LoadQueue.scala 152:68:@12703.4]
  wire  _T_14880; // @[LoadQueue.scala 151:92:@12705.4]
  wire  _T_14881; // @[LoadQueue.scala 152:41:@12706.4]
  wire  _T_14882; // @[LoadQueue.scala 153:30:@12707.4]
  wire  conflict_5_2; // @[LoadQueue.scala 152:68:@12708.4]
  wire  _T_14884; // @[LoadQueue.scala 151:92:@12710.4]
  wire  _T_14885; // @[LoadQueue.scala 152:41:@12711.4]
  wire  _T_14886; // @[LoadQueue.scala 153:30:@12712.4]
  wire  conflict_5_3; // @[LoadQueue.scala 152:68:@12713.4]
  wire  _T_14888; // @[LoadQueue.scala 151:92:@12715.4]
  wire  _T_14889; // @[LoadQueue.scala 152:41:@12716.4]
  wire  _T_14890; // @[LoadQueue.scala 153:30:@12717.4]
  wire  conflict_5_4; // @[LoadQueue.scala 152:68:@12718.4]
  wire  _T_14892; // @[LoadQueue.scala 151:92:@12720.4]
  wire  _T_14893; // @[LoadQueue.scala 152:41:@12721.4]
  wire  _T_14894; // @[LoadQueue.scala 153:30:@12722.4]
  wire  conflict_5_5; // @[LoadQueue.scala 152:68:@12723.4]
  wire  _T_14896; // @[LoadQueue.scala 151:92:@12725.4]
  wire  _T_14897; // @[LoadQueue.scala 152:41:@12726.4]
  wire  _T_14898; // @[LoadQueue.scala 153:30:@12727.4]
  wire  conflict_5_6; // @[LoadQueue.scala 152:68:@12728.4]
  wire  _T_14900; // @[LoadQueue.scala 151:92:@12730.4]
  wire  _T_14901; // @[LoadQueue.scala 152:41:@12731.4]
  wire  _T_14902; // @[LoadQueue.scala 153:30:@12732.4]
  wire  conflict_5_7; // @[LoadQueue.scala 152:68:@12733.4]
  wire  _T_14904; // @[LoadQueue.scala 151:92:@12735.4]
  wire  _T_14905; // @[LoadQueue.scala 152:41:@12736.4]
  wire  _T_14906; // @[LoadQueue.scala 153:30:@12737.4]
  wire  conflict_5_8; // @[LoadQueue.scala 152:68:@12738.4]
  wire  _T_14908; // @[LoadQueue.scala 151:92:@12740.4]
  wire  _T_14909; // @[LoadQueue.scala 152:41:@12741.4]
  wire  _T_14910; // @[LoadQueue.scala 153:30:@12742.4]
  wire  conflict_5_9; // @[LoadQueue.scala 152:68:@12743.4]
  wire  _T_14912; // @[LoadQueue.scala 151:92:@12745.4]
  wire  _T_14913; // @[LoadQueue.scala 152:41:@12746.4]
  wire  _T_14914; // @[LoadQueue.scala 153:30:@12747.4]
  wire  conflict_5_10; // @[LoadQueue.scala 152:68:@12748.4]
  wire  _T_14916; // @[LoadQueue.scala 151:92:@12750.4]
  wire  _T_14917; // @[LoadQueue.scala 152:41:@12751.4]
  wire  _T_14918; // @[LoadQueue.scala 153:30:@12752.4]
  wire  conflict_5_11; // @[LoadQueue.scala 152:68:@12753.4]
  wire  _T_14920; // @[LoadQueue.scala 151:92:@12755.4]
  wire  _T_14921; // @[LoadQueue.scala 152:41:@12756.4]
  wire  _T_14922; // @[LoadQueue.scala 153:30:@12757.4]
  wire  conflict_5_12; // @[LoadQueue.scala 152:68:@12758.4]
  wire  _T_14924; // @[LoadQueue.scala 151:92:@12760.4]
  wire  _T_14925; // @[LoadQueue.scala 152:41:@12761.4]
  wire  _T_14926; // @[LoadQueue.scala 153:30:@12762.4]
  wire  conflict_5_13; // @[LoadQueue.scala 152:68:@12763.4]
  wire  _T_14928; // @[LoadQueue.scala 151:92:@12765.4]
  wire  _T_14929; // @[LoadQueue.scala 152:41:@12766.4]
  wire  _T_14930; // @[LoadQueue.scala 153:30:@12767.4]
  wire  conflict_5_14; // @[LoadQueue.scala 152:68:@12768.4]
  wire  _T_14932; // @[LoadQueue.scala 151:92:@12770.4]
  wire  _T_14933; // @[LoadQueue.scala 152:41:@12771.4]
  wire  _T_14934; // @[LoadQueue.scala 153:30:@12772.4]
  wire  conflict_5_15; // @[LoadQueue.scala 152:68:@12773.4]
  wire  _T_14936; // @[LoadQueue.scala 151:92:@12775.4]
  wire  _T_14937; // @[LoadQueue.scala 152:41:@12776.4]
  wire  _T_14938; // @[LoadQueue.scala 153:30:@12777.4]
  wire  conflict_6_0; // @[LoadQueue.scala 152:68:@12778.4]
  wire  _T_14940; // @[LoadQueue.scala 151:92:@12780.4]
  wire  _T_14941; // @[LoadQueue.scala 152:41:@12781.4]
  wire  _T_14942; // @[LoadQueue.scala 153:30:@12782.4]
  wire  conflict_6_1; // @[LoadQueue.scala 152:68:@12783.4]
  wire  _T_14944; // @[LoadQueue.scala 151:92:@12785.4]
  wire  _T_14945; // @[LoadQueue.scala 152:41:@12786.4]
  wire  _T_14946; // @[LoadQueue.scala 153:30:@12787.4]
  wire  conflict_6_2; // @[LoadQueue.scala 152:68:@12788.4]
  wire  _T_14948; // @[LoadQueue.scala 151:92:@12790.4]
  wire  _T_14949; // @[LoadQueue.scala 152:41:@12791.4]
  wire  _T_14950; // @[LoadQueue.scala 153:30:@12792.4]
  wire  conflict_6_3; // @[LoadQueue.scala 152:68:@12793.4]
  wire  _T_14952; // @[LoadQueue.scala 151:92:@12795.4]
  wire  _T_14953; // @[LoadQueue.scala 152:41:@12796.4]
  wire  _T_14954; // @[LoadQueue.scala 153:30:@12797.4]
  wire  conflict_6_4; // @[LoadQueue.scala 152:68:@12798.4]
  wire  _T_14956; // @[LoadQueue.scala 151:92:@12800.4]
  wire  _T_14957; // @[LoadQueue.scala 152:41:@12801.4]
  wire  _T_14958; // @[LoadQueue.scala 153:30:@12802.4]
  wire  conflict_6_5; // @[LoadQueue.scala 152:68:@12803.4]
  wire  _T_14960; // @[LoadQueue.scala 151:92:@12805.4]
  wire  _T_14961; // @[LoadQueue.scala 152:41:@12806.4]
  wire  _T_14962; // @[LoadQueue.scala 153:30:@12807.4]
  wire  conflict_6_6; // @[LoadQueue.scala 152:68:@12808.4]
  wire  _T_14964; // @[LoadQueue.scala 151:92:@12810.4]
  wire  _T_14965; // @[LoadQueue.scala 152:41:@12811.4]
  wire  _T_14966; // @[LoadQueue.scala 153:30:@12812.4]
  wire  conflict_6_7; // @[LoadQueue.scala 152:68:@12813.4]
  wire  _T_14968; // @[LoadQueue.scala 151:92:@12815.4]
  wire  _T_14969; // @[LoadQueue.scala 152:41:@12816.4]
  wire  _T_14970; // @[LoadQueue.scala 153:30:@12817.4]
  wire  conflict_6_8; // @[LoadQueue.scala 152:68:@12818.4]
  wire  _T_14972; // @[LoadQueue.scala 151:92:@12820.4]
  wire  _T_14973; // @[LoadQueue.scala 152:41:@12821.4]
  wire  _T_14974; // @[LoadQueue.scala 153:30:@12822.4]
  wire  conflict_6_9; // @[LoadQueue.scala 152:68:@12823.4]
  wire  _T_14976; // @[LoadQueue.scala 151:92:@12825.4]
  wire  _T_14977; // @[LoadQueue.scala 152:41:@12826.4]
  wire  _T_14978; // @[LoadQueue.scala 153:30:@12827.4]
  wire  conflict_6_10; // @[LoadQueue.scala 152:68:@12828.4]
  wire  _T_14980; // @[LoadQueue.scala 151:92:@12830.4]
  wire  _T_14981; // @[LoadQueue.scala 152:41:@12831.4]
  wire  _T_14982; // @[LoadQueue.scala 153:30:@12832.4]
  wire  conflict_6_11; // @[LoadQueue.scala 152:68:@12833.4]
  wire  _T_14984; // @[LoadQueue.scala 151:92:@12835.4]
  wire  _T_14985; // @[LoadQueue.scala 152:41:@12836.4]
  wire  _T_14986; // @[LoadQueue.scala 153:30:@12837.4]
  wire  conflict_6_12; // @[LoadQueue.scala 152:68:@12838.4]
  wire  _T_14988; // @[LoadQueue.scala 151:92:@12840.4]
  wire  _T_14989; // @[LoadQueue.scala 152:41:@12841.4]
  wire  _T_14990; // @[LoadQueue.scala 153:30:@12842.4]
  wire  conflict_6_13; // @[LoadQueue.scala 152:68:@12843.4]
  wire  _T_14992; // @[LoadQueue.scala 151:92:@12845.4]
  wire  _T_14993; // @[LoadQueue.scala 152:41:@12846.4]
  wire  _T_14994; // @[LoadQueue.scala 153:30:@12847.4]
  wire  conflict_6_14; // @[LoadQueue.scala 152:68:@12848.4]
  wire  _T_14996; // @[LoadQueue.scala 151:92:@12850.4]
  wire  _T_14997; // @[LoadQueue.scala 152:41:@12851.4]
  wire  _T_14998; // @[LoadQueue.scala 153:30:@12852.4]
  wire  conflict_6_15; // @[LoadQueue.scala 152:68:@12853.4]
  wire  _T_15000; // @[LoadQueue.scala 151:92:@12855.4]
  wire  _T_15001; // @[LoadQueue.scala 152:41:@12856.4]
  wire  _T_15002; // @[LoadQueue.scala 153:30:@12857.4]
  wire  conflict_7_0; // @[LoadQueue.scala 152:68:@12858.4]
  wire  _T_15004; // @[LoadQueue.scala 151:92:@12860.4]
  wire  _T_15005; // @[LoadQueue.scala 152:41:@12861.4]
  wire  _T_15006; // @[LoadQueue.scala 153:30:@12862.4]
  wire  conflict_7_1; // @[LoadQueue.scala 152:68:@12863.4]
  wire  _T_15008; // @[LoadQueue.scala 151:92:@12865.4]
  wire  _T_15009; // @[LoadQueue.scala 152:41:@12866.4]
  wire  _T_15010; // @[LoadQueue.scala 153:30:@12867.4]
  wire  conflict_7_2; // @[LoadQueue.scala 152:68:@12868.4]
  wire  _T_15012; // @[LoadQueue.scala 151:92:@12870.4]
  wire  _T_15013; // @[LoadQueue.scala 152:41:@12871.4]
  wire  _T_15014; // @[LoadQueue.scala 153:30:@12872.4]
  wire  conflict_7_3; // @[LoadQueue.scala 152:68:@12873.4]
  wire  _T_15016; // @[LoadQueue.scala 151:92:@12875.4]
  wire  _T_15017; // @[LoadQueue.scala 152:41:@12876.4]
  wire  _T_15018; // @[LoadQueue.scala 153:30:@12877.4]
  wire  conflict_7_4; // @[LoadQueue.scala 152:68:@12878.4]
  wire  _T_15020; // @[LoadQueue.scala 151:92:@12880.4]
  wire  _T_15021; // @[LoadQueue.scala 152:41:@12881.4]
  wire  _T_15022; // @[LoadQueue.scala 153:30:@12882.4]
  wire  conflict_7_5; // @[LoadQueue.scala 152:68:@12883.4]
  wire  _T_15024; // @[LoadQueue.scala 151:92:@12885.4]
  wire  _T_15025; // @[LoadQueue.scala 152:41:@12886.4]
  wire  _T_15026; // @[LoadQueue.scala 153:30:@12887.4]
  wire  conflict_7_6; // @[LoadQueue.scala 152:68:@12888.4]
  wire  _T_15028; // @[LoadQueue.scala 151:92:@12890.4]
  wire  _T_15029; // @[LoadQueue.scala 152:41:@12891.4]
  wire  _T_15030; // @[LoadQueue.scala 153:30:@12892.4]
  wire  conflict_7_7; // @[LoadQueue.scala 152:68:@12893.4]
  wire  _T_15032; // @[LoadQueue.scala 151:92:@12895.4]
  wire  _T_15033; // @[LoadQueue.scala 152:41:@12896.4]
  wire  _T_15034; // @[LoadQueue.scala 153:30:@12897.4]
  wire  conflict_7_8; // @[LoadQueue.scala 152:68:@12898.4]
  wire  _T_15036; // @[LoadQueue.scala 151:92:@12900.4]
  wire  _T_15037; // @[LoadQueue.scala 152:41:@12901.4]
  wire  _T_15038; // @[LoadQueue.scala 153:30:@12902.4]
  wire  conflict_7_9; // @[LoadQueue.scala 152:68:@12903.4]
  wire  _T_15040; // @[LoadQueue.scala 151:92:@12905.4]
  wire  _T_15041; // @[LoadQueue.scala 152:41:@12906.4]
  wire  _T_15042; // @[LoadQueue.scala 153:30:@12907.4]
  wire  conflict_7_10; // @[LoadQueue.scala 152:68:@12908.4]
  wire  _T_15044; // @[LoadQueue.scala 151:92:@12910.4]
  wire  _T_15045; // @[LoadQueue.scala 152:41:@12911.4]
  wire  _T_15046; // @[LoadQueue.scala 153:30:@12912.4]
  wire  conflict_7_11; // @[LoadQueue.scala 152:68:@12913.4]
  wire  _T_15048; // @[LoadQueue.scala 151:92:@12915.4]
  wire  _T_15049; // @[LoadQueue.scala 152:41:@12916.4]
  wire  _T_15050; // @[LoadQueue.scala 153:30:@12917.4]
  wire  conflict_7_12; // @[LoadQueue.scala 152:68:@12918.4]
  wire  _T_15052; // @[LoadQueue.scala 151:92:@12920.4]
  wire  _T_15053; // @[LoadQueue.scala 152:41:@12921.4]
  wire  _T_15054; // @[LoadQueue.scala 153:30:@12922.4]
  wire  conflict_7_13; // @[LoadQueue.scala 152:68:@12923.4]
  wire  _T_15056; // @[LoadQueue.scala 151:92:@12925.4]
  wire  _T_15057; // @[LoadQueue.scala 152:41:@12926.4]
  wire  _T_15058; // @[LoadQueue.scala 153:30:@12927.4]
  wire  conflict_7_14; // @[LoadQueue.scala 152:68:@12928.4]
  wire  _T_15060; // @[LoadQueue.scala 151:92:@12930.4]
  wire  _T_15061; // @[LoadQueue.scala 152:41:@12931.4]
  wire  _T_15062; // @[LoadQueue.scala 153:30:@12932.4]
  wire  conflict_7_15; // @[LoadQueue.scala 152:68:@12933.4]
  wire  _T_15064; // @[LoadQueue.scala 151:92:@12935.4]
  wire  _T_15065; // @[LoadQueue.scala 152:41:@12936.4]
  wire  _T_15066; // @[LoadQueue.scala 153:30:@12937.4]
  wire  conflict_8_0; // @[LoadQueue.scala 152:68:@12938.4]
  wire  _T_15068; // @[LoadQueue.scala 151:92:@12940.4]
  wire  _T_15069; // @[LoadQueue.scala 152:41:@12941.4]
  wire  _T_15070; // @[LoadQueue.scala 153:30:@12942.4]
  wire  conflict_8_1; // @[LoadQueue.scala 152:68:@12943.4]
  wire  _T_15072; // @[LoadQueue.scala 151:92:@12945.4]
  wire  _T_15073; // @[LoadQueue.scala 152:41:@12946.4]
  wire  _T_15074; // @[LoadQueue.scala 153:30:@12947.4]
  wire  conflict_8_2; // @[LoadQueue.scala 152:68:@12948.4]
  wire  _T_15076; // @[LoadQueue.scala 151:92:@12950.4]
  wire  _T_15077; // @[LoadQueue.scala 152:41:@12951.4]
  wire  _T_15078; // @[LoadQueue.scala 153:30:@12952.4]
  wire  conflict_8_3; // @[LoadQueue.scala 152:68:@12953.4]
  wire  _T_15080; // @[LoadQueue.scala 151:92:@12955.4]
  wire  _T_15081; // @[LoadQueue.scala 152:41:@12956.4]
  wire  _T_15082; // @[LoadQueue.scala 153:30:@12957.4]
  wire  conflict_8_4; // @[LoadQueue.scala 152:68:@12958.4]
  wire  _T_15084; // @[LoadQueue.scala 151:92:@12960.4]
  wire  _T_15085; // @[LoadQueue.scala 152:41:@12961.4]
  wire  _T_15086; // @[LoadQueue.scala 153:30:@12962.4]
  wire  conflict_8_5; // @[LoadQueue.scala 152:68:@12963.4]
  wire  _T_15088; // @[LoadQueue.scala 151:92:@12965.4]
  wire  _T_15089; // @[LoadQueue.scala 152:41:@12966.4]
  wire  _T_15090; // @[LoadQueue.scala 153:30:@12967.4]
  wire  conflict_8_6; // @[LoadQueue.scala 152:68:@12968.4]
  wire  _T_15092; // @[LoadQueue.scala 151:92:@12970.4]
  wire  _T_15093; // @[LoadQueue.scala 152:41:@12971.4]
  wire  _T_15094; // @[LoadQueue.scala 153:30:@12972.4]
  wire  conflict_8_7; // @[LoadQueue.scala 152:68:@12973.4]
  wire  _T_15096; // @[LoadQueue.scala 151:92:@12975.4]
  wire  _T_15097; // @[LoadQueue.scala 152:41:@12976.4]
  wire  _T_15098; // @[LoadQueue.scala 153:30:@12977.4]
  wire  conflict_8_8; // @[LoadQueue.scala 152:68:@12978.4]
  wire  _T_15100; // @[LoadQueue.scala 151:92:@12980.4]
  wire  _T_15101; // @[LoadQueue.scala 152:41:@12981.4]
  wire  _T_15102; // @[LoadQueue.scala 153:30:@12982.4]
  wire  conflict_8_9; // @[LoadQueue.scala 152:68:@12983.4]
  wire  _T_15104; // @[LoadQueue.scala 151:92:@12985.4]
  wire  _T_15105; // @[LoadQueue.scala 152:41:@12986.4]
  wire  _T_15106; // @[LoadQueue.scala 153:30:@12987.4]
  wire  conflict_8_10; // @[LoadQueue.scala 152:68:@12988.4]
  wire  _T_15108; // @[LoadQueue.scala 151:92:@12990.4]
  wire  _T_15109; // @[LoadQueue.scala 152:41:@12991.4]
  wire  _T_15110; // @[LoadQueue.scala 153:30:@12992.4]
  wire  conflict_8_11; // @[LoadQueue.scala 152:68:@12993.4]
  wire  _T_15112; // @[LoadQueue.scala 151:92:@12995.4]
  wire  _T_15113; // @[LoadQueue.scala 152:41:@12996.4]
  wire  _T_15114; // @[LoadQueue.scala 153:30:@12997.4]
  wire  conflict_8_12; // @[LoadQueue.scala 152:68:@12998.4]
  wire  _T_15116; // @[LoadQueue.scala 151:92:@13000.4]
  wire  _T_15117; // @[LoadQueue.scala 152:41:@13001.4]
  wire  _T_15118; // @[LoadQueue.scala 153:30:@13002.4]
  wire  conflict_8_13; // @[LoadQueue.scala 152:68:@13003.4]
  wire  _T_15120; // @[LoadQueue.scala 151:92:@13005.4]
  wire  _T_15121; // @[LoadQueue.scala 152:41:@13006.4]
  wire  _T_15122; // @[LoadQueue.scala 153:30:@13007.4]
  wire  conflict_8_14; // @[LoadQueue.scala 152:68:@13008.4]
  wire  _T_15124; // @[LoadQueue.scala 151:92:@13010.4]
  wire  _T_15125; // @[LoadQueue.scala 152:41:@13011.4]
  wire  _T_15126; // @[LoadQueue.scala 153:30:@13012.4]
  wire  conflict_8_15; // @[LoadQueue.scala 152:68:@13013.4]
  wire  _T_15128; // @[LoadQueue.scala 151:92:@13015.4]
  wire  _T_15129; // @[LoadQueue.scala 152:41:@13016.4]
  wire  _T_15130; // @[LoadQueue.scala 153:30:@13017.4]
  wire  conflict_9_0; // @[LoadQueue.scala 152:68:@13018.4]
  wire  _T_15132; // @[LoadQueue.scala 151:92:@13020.4]
  wire  _T_15133; // @[LoadQueue.scala 152:41:@13021.4]
  wire  _T_15134; // @[LoadQueue.scala 153:30:@13022.4]
  wire  conflict_9_1; // @[LoadQueue.scala 152:68:@13023.4]
  wire  _T_15136; // @[LoadQueue.scala 151:92:@13025.4]
  wire  _T_15137; // @[LoadQueue.scala 152:41:@13026.4]
  wire  _T_15138; // @[LoadQueue.scala 153:30:@13027.4]
  wire  conflict_9_2; // @[LoadQueue.scala 152:68:@13028.4]
  wire  _T_15140; // @[LoadQueue.scala 151:92:@13030.4]
  wire  _T_15141; // @[LoadQueue.scala 152:41:@13031.4]
  wire  _T_15142; // @[LoadQueue.scala 153:30:@13032.4]
  wire  conflict_9_3; // @[LoadQueue.scala 152:68:@13033.4]
  wire  _T_15144; // @[LoadQueue.scala 151:92:@13035.4]
  wire  _T_15145; // @[LoadQueue.scala 152:41:@13036.4]
  wire  _T_15146; // @[LoadQueue.scala 153:30:@13037.4]
  wire  conflict_9_4; // @[LoadQueue.scala 152:68:@13038.4]
  wire  _T_15148; // @[LoadQueue.scala 151:92:@13040.4]
  wire  _T_15149; // @[LoadQueue.scala 152:41:@13041.4]
  wire  _T_15150; // @[LoadQueue.scala 153:30:@13042.4]
  wire  conflict_9_5; // @[LoadQueue.scala 152:68:@13043.4]
  wire  _T_15152; // @[LoadQueue.scala 151:92:@13045.4]
  wire  _T_15153; // @[LoadQueue.scala 152:41:@13046.4]
  wire  _T_15154; // @[LoadQueue.scala 153:30:@13047.4]
  wire  conflict_9_6; // @[LoadQueue.scala 152:68:@13048.4]
  wire  _T_15156; // @[LoadQueue.scala 151:92:@13050.4]
  wire  _T_15157; // @[LoadQueue.scala 152:41:@13051.4]
  wire  _T_15158; // @[LoadQueue.scala 153:30:@13052.4]
  wire  conflict_9_7; // @[LoadQueue.scala 152:68:@13053.4]
  wire  _T_15160; // @[LoadQueue.scala 151:92:@13055.4]
  wire  _T_15161; // @[LoadQueue.scala 152:41:@13056.4]
  wire  _T_15162; // @[LoadQueue.scala 153:30:@13057.4]
  wire  conflict_9_8; // @[LoadQueue.scala 152:68:@13058.4]
  wire  _T_15164; // @[LoadQueue.scala 151:92:@13060.4]
  wire  _T_15165; // @[LoadQueue.scala 152:41:@13061.4]
  wire  _T_15166; // @[LoadQueue.scala 153:30:@13062.4]
  wire  conflict_9_9; // @[LoadQueue.scala 152:68:@13063.4]
  wire  _T_15168; // @[LoadQueue.scala 151:92:@13065.4]
  wire  _T_15169; // @[LoadQueue.scala 152:41:@13066.4]
  wire  _T_15170; // @[LoadQueue.scala 153:30:@13067.4]
  wire  conflict_9_10; // @[LoadQueue.scala 152:68:@13068.4]
  wire  _T_15172; // @[LoadQueue.scala 151:92:@13070.4]
  wire  _T_15173; // @[LoadQueue.scala 152:41:@13071.4]
  wire  _T_15174; // @[LoadQueue.scala 153:30:@13072.4]
  wire  conflict_9_11; // @[LoadQueue.scala 152:68:@13073.4]
  wire  _T_15176; // @[LoadQueue.scala 151:92:@13075.4]
  wire  _T_15177; // @[LoadQueue.scala 152:41:@13076.4]
  wire  _T_15178; // @[LoadQueue.scala 153:30:@13077.4]
  wire  conflict_9_12; // @[LoadQueue.scala 152:68:@13078.4]
  wire  _T_15180; // @[LoadQueue.scala 151:92:@13080.4]
  wire  _T_15181; // @[LoadQueue.scala 152:41:@13081.4]
  wire  _T_15182; // @[LoadQueue.scala 153:30:@13082.4]
  wire  conflict_9_13; // @[LoadQueue.scala 152:68:@13083.4]
  wire  _T_15184; // @[LoadQueue.scala 151:92:@13085.4]
  wire  _T_15185; // @[LoadQueue.scala 152:41:@13086.4]
  wire  _T_15186; // @[LoadQueue.scala 153:30:@13087.4]
  wire  conflict_9_14; // @[LoadQueue.scala 152:68:@13088.4]
  wire  _T_15188; // @[LoadQueue.scala 151:92:@13090.4]
  wire  _T_15189; // @[LoadQueue.scala 152:41:@13091.4]
  wire  _T_15190; // @[LoadQueue.scala 153:30:@13092.4]
  wire  conflict_9_15; // @[LoadQueue.scala 152:68:@13093.4]
  wire  _T_15192; // @[LoadQueue.scala 151:92:@13095.4]
  wire  _T_15193; // @[LoadQueue.scala 152:41:@13096.4]
  wire  _T_15194; // @[LoadQueue.scala 153:30:@13097.4]
  wire  conflict_10_0; // @[LoadQueue.scala 152:68:@13098.4]
  wire  _T_15196; // @[LoadQueue.scala 151:92:@13100.4]
  wire  _T_15197; // @[LoadQueue.scala 152:41:@13101.4]
  wire  _T_15198; // @[LoadQueue.scala 153:30:@13102.4]
  wire  conflict_10_1; // @[LoadQueue.scala 152:68:@13103.4]
  wire  _T_15200; // @[LoadQueue.scala 151:92:@13105.4]
  wire  _T_15201; // @[LoadQueue.scala 152:41:@13106.4]
  wire  _T_15202; // @[LoadQueue.scala 153:30:@13107.4]
  wire  conflict_10_2; // @[LoadQueue.scala 152:68:@13108.4]
  wire  _T_15204; // @[LoadQueue.scala 151:92:@13110.4]
  wire  _T_15205; // @[LoadQueue.scala 152:41:@13111.4]
  wire  _T_15206; // @[LoadQueue.scala 153:30:@13112.4]
  wire  conflict_10_3; // @[LoadQueue.scala 152:68:@13113.4]
  wire  _T_15208; // @[LoadQueue.scala 151:92:@13115.4]
  wire  _T_15209; // @[LoadQueue.scala 152:41:@13116.4]
  wire  _T_15210; // @[LoadQueue.scala 153:30:@13117.4]
  wire  conflict_10_4; // @[LoadQueue.scala 152:68:@13118.4]
  wire  _T_15212; // @[LoadQueue.scala 151:92:@13120.4]
  wire  _T_15213; // @[LoadQueue.scala 152:41:@13121.4]
  wire  _T_15214; // @[LoadQueue.scala 153:30:@13122.4]
  wire  conflict_10_5; // @[LoadQueue.scala 152:68:@13123.4]
  wire  _T_15216; // @[LoadQueue.scala 151:92:@13125.4]
  wire  _T_15217; // @[LoadQueue.scala 152:41:@13126.4]
  wire  _T_15218; // @[LoadQueue.scala 153:30:@13127.4]
  wire  conflict_10_6; // @[LoadQueue.scala 152:68:@13128.4]
  wire  _T_15220; // @[LoadQueue.scala 151:92:@13130.4]
  wire  _T_15221; // @[LoadQueue.scala 152:41:@13131.4]
  wire  _T_15222; // @[LoadQueue.scala 153:30:@13132.4]
  wire  conflict_10_7; // @[LoadQueue.scala 152:68:@13133.4]
  wire  _T_15224; // @[LoadQueue.scala 151:92:@13135.4]
  wire  _T_15225; // @[LoadQueue.scala 152:41:@13136.4]
  wire  _T_15226; // @[LoadQueue.scala 153:30:@13137.4]
  wire  conflict_10_8; // @[LoadQueue.scala 152:68:@13138.4]
  wire  _T_15228; // @[LoadQueue.scala 151:92:@13140.4]
  wire  _T_15229; // @[LoadQueue.scala 152:41:@13141.4]
  wire  _T_15230; // @[LoadQueue.scala 153:30:@13142.4]
  wire  conflict_10_9; // @[LoadQueue.scala 152:68:@13143.4]
  wire  _T_15232; // @[LoadQueue.scala 151:92:@13145.4]
  wire  _T_15233; // @[LoadQueue.scala 152:41:@13146.4]
  wire  _T_15234; // @[LoadQueue.scala 153:30:@13147.4]
  wire  conflict_10_10; // @[LoadQueue.scala 152:68:@13148.4]
  wire  _T_15236; // @[LoadQueue.scala 151:92:@13150.4]
  wire  _T_15237; // @[LoadQueue.scala 152:41:@13151.4]
  wire  _T_15238; // @[LoadQueue.scala 153:30:@13152.4]
  wire  conflict_10_11; // @[LoadQueue.scala 152:68:@13153.4]
  wire  _T_15240; // @[LoadQueue.scala 151:92:@13155.4]
  wire  _T_15241; // @[LoadQueue.scala 152:41:@13156.4]
  wire  _T_15242; // @[LoadQueue.scala 153:30:@13157.4]
  wire  conflict_10_12; // @[LoadQueue.scala 152:68:@13158.4]
  wire  _T_15244; // @[LoadQueue.scala 151:92:@13160.4]
  wire  _T_15245; // @[LoadQueue.scala 152:41:@13161.4]
  wire  _T_15246; // @[LoadQueue.scala 153:30:@13162.4]
  wire  conflict_10_13; // @[LoadQueue.scala 152:68:@13163.4]
  wire  _T_15248; // @[LoadQueue.scala 151:92:@13165.4]
  wire  _T_15249; // @[LoadQueue.scala 152:41:@13166.4]
  wire  _T_15250; // @[LoadQueue.scala 153:30:@13167.4]
  wire  conflict_10_14; // @[LoadQueue.scala 152:68:@13168.4]
  wire  _T_15252; // @[LoadQueue.scala 151:92:@13170.4]
  wire  _T_15253; // @[LoadQueue.scala 152:41:@13171.4]
  wire  _T_15254; // @[LoadQueue.scala 153:30:@13172.4]
  wire  conflict_10_15; // @[LoadQueue.scala 152:68:@13173.4]
  wire  _T_15256; // @[LoadQueue.scala 151:92:@13175.4]
  wire  _T_15257; // @[LoadQueue.scala 152:41:@13176.4]
  wire  _T_15258; // @[LoadQueue.scala 153:30:@13177.4]
  wire  conflict_11_0; // @[LoadQueue.scala 152:68:@13178.4]
  wire  _T_15260; // @[LoadQueue.scala 151:92:@13180.4]
  wire  _T_15261; // @[LoadQueue.scala 152:41:@13181.4]
  wire  _T_15262; // @[LoadQueue.scala 153:30:@13182.4]
  wire  conflict_11_1; // @[LoadQueue.scala 152:68:@13183.4]
  wire  _T_15264; // @[LoadQueue.scala 151:92:@13185.4]
  wire  _T_15265; // @[LoadQueue.scala 152:41:@13186.4]
  wire  _T_15266; // @[LoadQueue.scala 153:30:@13187.4]
  wire  conflict_11_2; // @[LoadQueue.scala 152:68:@13188.4]
  wire  _T_15268; // @[LoadQueue.scala 151:92:@13190.4]
  wire  _T_15269; // @[LoadQueue.scala 152:41:@13191.4]
  wire  _T_15270; // @[LoadQueue.scala 153:30:@13192.4]
  wire  conflict_11_3; // @[LoadQueue.scala 152:68:@13193.4]
  wire  _T_15272; // @[LoadQueue.scala 151:92:@13195.4]
  wire  _T_15273; // @[LoadQueue.scala 152:41:@13196.4]
  wire  _T_15274; // @[LoadQueue.scala 153:30:@13197.4]
  wire  conflict_11_4; // @[LoadQueue.scala 152:68:@13198.4]
  wire  _T_15276; // @[LoadQueue.scala 151:92:@13200.4]
  wire  _T_15277; // @[LoadQueue.scala 152:41:@13201.4]
  wire  _T_15278; // @[LoadQueue.scala 153:30:@13202.4]
  wire  conflict_11_5; // @[LoadQueue.scala 152:68:@13203.4]
  wire  _T_15280; // @[LoadQueue.scala 151:92:@13205.4]
  wire  _T_15281; // @[LoadQueue.scala 152:41:@13206.4]
  wire  _T_15282; // @[LoadQueue.scala 153:30:@13207.4]
  wire  conflict_11_6; // @[LoadQueue.scala 152:68:@13208.4]
  wire  _T_15284; // @[LoadQueue.scala 151:92:@13210.4]
  wire  _T_15285; // @[LoadQueue.scala 152:41:@13211.4]
  wire  _T_15286; // @[LoadQueue.scala 153:30:@13212.4]
  wire  conflict_11_7; // @[LoadQueue.scala 152:68:@13213.4]
  wire  _T_15288; // @[LoadQueue.scala 151:92:@13215.4]
  wire  _T_15289; // @[LoadQueue.scala 152:41:@13216.4]
  wire  _T_15290; // @[LoadQueue.scala 153:30:@13217.4]
  wire  conflict_11_8; // @[LoadQueue.scala 152:68:@13218.4]
  wire  _T_15292; // @[LoadQueue.scala 151:92:@13220.4]
  wire  _T_15293; // @[LoadQueue.scala 152:41:@13221.4]
  wire  _T_15294; // @[LoadQueue.scala 153:30:@13222.4]
  wire  conflict_11_9; // @[LoadQueue.scala 152:68:@13223.4]
  wire  _T_15296; // @[LoadQueue.scala 151:92:@13225.4]
  wire  _T_15297; // @[LoadQueue.scala 152:41:@13226.4]
  wire  _T_15298; // @[LoadQueue.scala 153:30:@13227.4]
  wire  conflict_11_10; // @[LoadQueue.scala 152:68:@13228.4]
  wire  _T_15300; // @[LoadQueue.scala 151:92:@13230.4]
  wire  _T_15301; // @[LoadQueue.scala 152:41:@13231.4]
  wire  _T_15302; // @[LoadQueue.scala 153:30:@13232.4]
  wire  conflict_11_11; // @[LoadQueue.scala 152:68:@13233.4]
  wire  _T_15304; // @[LoadQueue.scala 151:92:@13235.4]
  wire  _T_15305; // @[LoadQueue.scala 152:41:@13236.4]
  wire  _T_15306; // @[LoadQueue.scala 153:30:@13237.4]
  wire  conflict_11_12; // @[LoadQueue.scala 152:68:@13238.4]
  wire  _T_15308; // @[LoadQueue.scala 151:92:@13240.4]
  wire  _T_15309; // @[LoadQueue.scala 152:41:@13241.4]
  wire  _T_15310; // @[LoadQueue.scala 153:30:@13242.4]
  wire  conflict_11_13; // @[LoadQueue.scala 152:68:@13243.4]
  wire  _T_15312; // @[LoadQueue.scala 151:92:@13245.4]
  wire  _T_15313; // @[LoadQueue.scala 152:41:@13246.4]
  wire  _T_15314; // @[LoadQueue.scala 153:30:@13247.4]
  wire  conflict_11_14; // @[LoadQueue.scala 152:68:@13248.4]
  wire  _T_15316; // @[LoadQueue.scala 151:92:@13250.4]
  wire  _T_15317; // @[LoadQueue.scala 152:41:@13251.4]
  wire  _T_15318; // @[LoadQueue.scala 153:30:@13252.4]
  wire  conflict_11_15; // @[LoadQueue.scala 152:68:@13253.4]
  wire  _T_15320; // @[LoadQueue.scala 151:92:@13255.4]
  wire  _T_15321; // @[LoadQueue.scala 152:41:@13256.4]
  wire  _T_15322; // @[LoadQueue.scala 153:30:@13257.4]
  wire  conflict_12_0; // @[LoadQueue.scala 152:68:@13258.4]
  wire  _T_15324; // @[LoadQueue.scala 151:92:@13260.4]
  wire  _T_15325; // @[LoadQueue.scala 152:41:@13261.4]
  wire  _T_15326; // @[LoadQueue.scala 153:30:@13262.4]
  wire  conflict_12_1; // @[LoadQueue.scala 152:68:@13263.4]
  wire  _T_15328; // @[LoadQueue.scala 151:92:@13265.4]
  wire  _T_15329; // @[LoadQueue.scala 152:41:@13266.4]
  wire  _T_15330; // @[LoadQueue.scala 153:30:@13267.4]
  wire  conflict_12_2; // @[LoadQueue.scala 152:68:@13268.4]
  wire  _T_15332; // @[LoadQueue.scala 151:92:@13270.4]
  wire  _T_15333; // @[LoadQueue.scala 152:41:@13271.4]
  wire  _T_15334; // @[LoadQueue.scala 153:30:@13272.4]
  wire  conflict_12_3; // @[LoadQueue.scala 152:68:@13273.4]
  wire  _T_15336; // @[LoadQueue.scala 151:92:@13275.4]
  wire  _T_15337; // @[LoadQueue.scala 152:41:@13276.4]
  wire  _T_15338; // @[LoadQueue.scala 153:30:@13277.4]
  wire  conflict_12_4; // @[LoadQueue.scala 152:68:@13278.4]
  wire  _T_15340; // @[LoadQueue.scala 151:92:@13280.4]
  wire  _T_15341; // @[LoadQueue.scala 152:41:@13281.4]
  wire  _T_15342; // @[LoadQueue.scala 153:30:@13282.4]
  wire  conflict_12_5; // @[LoadQueue.scala 152:68:@13283.4]
  wire  _T_15344; // @[LoadQueue.scala 151:92:@13285.4]
  wire  _T_15345; // @[LoadQueue.scala 152:41:@13286.4]
  wire  _T_15346; // @[LoadQueue.scala 153:30:@13287.4]
  wire  conflict_12_6; // @[LoadQueue.scala 152:68:@13288.4]
  wire  _T_15348; // @[LoadQueue.scala 151:92:@13290.4]
  wire  _T_15349; // @[LoadQueue.scala 152:41:@13291.4]
  wire  _T_15350; // @[LoadQueue.scala 153:30:@13292.4]
  wire  conflict_12_7; // @[LoadQueue.scala 152:68:@13293.4]
  wire  _T_15352; // @[LoadQueue.scala 151:92:@13295.4]
  wire  _T_15353; // @[LoadQueue.scala 152:41:@13296.4]
  wire  _T_15354; // @[LoadQueue.scala 153:30:@13297.4]
  wire  conflict_12_8; // @[LoadQueue.scala 152:68:@13298.4]
  wire  _T_15356; // @[LoadQueue.scala 151:92:@13300.4]
  wire  _T_15357; // @[LoadQueue.scala 152:41:@13301.4]
  wire  _T_15358; // @[LoadQueue.scala 153:30:@13302.4]
  wire  conflict_12_9; // @[LoadQueue.scala 152:68:@13303.4]
  wire  _T_15360; // @[LoadQueue.scala 151:92:@13305.4]
  wire  _T_15361; // @[LoadQueue.scala 152:41:@13306.4]
  wire  _T_15362; // @[LoadQueue.scala 153:30:@13307.4]
  wire  conflict_12_10; // @[LoadQueue.scala 152:68:@13308.4]
  wire  _T_15364; // @[LoadQueue.scala 151:92:@13310.4]
  wire  _T_15365; // @[LoadQueue.scala 152:41:@13311.4]
  wire  _T_15366; // @[LoadQueue.scala 153:30:@13312.4]
  wire  conflict_12_11; // @[LoadQueue.scala 152:68:@13313.4]
  wire  _T_15368; // @[LoadQueue.scala 151:92:@13315.4]
  wire  _T_15369; // @[LoadQueue.scala 152:41:@13316.4]
  wire  _T_15370; // @[LoadQueue.scala 153:30:@13317.4]
  wire  conflict_12_12; // @[LoadQueue.scala 152:68:@13318.4]
  wire  _T_15372; // @[LoadQueue.scala 151:92:@13320.4]
  wire  _T_15373; // @[LoadQueue.scala 152:41:@13321.4]
  wire  _T_15374; // @[LoadQueue.scala 153:30:@13322.4]
  wire  conflict_12_13; // @[LoadQueue.scala 152:68:@13323.4]
  wire  _T_15376; // @[LoadQueue.scala 151:92:@13325.4]
  wire  _T_15377; // @[LoadQueue.scala 152:41:@13326.4]
  wire  _T_15378; // @[LoadQueue.scala 153:30:@13327.4]
  wire  conflict_12_14; // @[LoadQueue.scala 152:68:@13328.4]
  wire  _T_15380; // @[LoadQueue.scala 151:92:@13330.4]
  wire  _T_15381; // @[LoadQueue.scala 152:41:@13331.4]
  wire  _T_15382; // @[LoadQueue.scala 153:30:@13332.4]
  wire  conflict_12_15; // @[LoadQueue.scala 152:68:@13333.4]
  wire  _T_15384; // @[LoadQueue.scala 151:92:@13335.4]
  wire  _T_15385; // @[LoadQueue.scala 152:41:@13336.4]
  wire  _T_15386; // @[LoadQueue.scala 153:30:@13337.4]
  wire  conflict_13_0; // @[LoadQueue.scala 152:68:@13338.4]
  wire  _T_15388; // @[LoadQueue.scala 151:92:@13340.4]
  wire  _T_15389; // @[LoadQueue.scala 152:41:@13341.4]
  wire  _T_15390; // @[LoadQueue.scala 153:30:@13342.4]
  wire  conflict_13_1; // @[LoadQueue.scala 152:68:@13343.4]
  wire  _T_15392; // @[LoadQueue.scala 151:92:@13345.4]
  wire  _T_15393; // @[LoadQueue.scala 152:41:@13346.4]
  wire  _T_15394; // @[LoadQueue.scala 153:30:@13347.4]
  wire  conflict_13_2; // @[LoadQueue.scala 152:68:@13348.4]
  wire  _T_15396; // @[LoadQueue.scala 151:92:@13350.4]
  wire  _T_15397; // @[LoadQueue.scala 152:41:@13351.4]
  wire  _T_15398; // @[LoadQueue.scala 153:30:@13352.4]
  wire  conflict_13_3; // @[LoadQueue.scala 152:68:@13353.4]
  wire  _T_15400; // @[LoadQueue.scala 151:92:@13355.4]
  wire  _T_15401; // @[LoadQueue.scala 152:41:@13356.4]
  wire  _T_15402; // @[LoadQueue.scala 153:30:@13357.4]
  wire  conflict_13_4; // @[LoadQueue.scala 152:68:@13358.4]
  wire  _T_15404; // @[LoadQueue.scala 151:92:@13360.4]
  wire  _T_15405; // @[LoadQueue.scala 152:41:@13361.4]
  wire  _T_15406; // @[LoadQueue.scala 153:30:@13362.4]
  wire  conflict_13_5; // @[LoadQueue.scala 152:68:@13363.4]
  wire  _T_15408; // @[LoadQueue.scala 151:92:@13365.4]
  wire  _T_15409; // @[LoadQueue.scala 152:41:@13366.4]
  wire  _T_15410; // @[LoadQueue.scala 153:30:@13367.4]
  wire  conflict_13_6; // @[LoadQueue.scala 152:68:@13368.4]
  wire  _T_15412; // @[LoadQueue.scala 151:92:@13370.4]
  wire  _T_15413; // @[LoadQueue.scala 152:41:@13371.4]
  wire  _T_15414; // @[LoadQueue.scala 153:30:@13372.4]
  wire  conflict_13_7; // @[LoadQueue.scala 152:68:@13373.4]
  wire  _T_15416; // @[LoadQueue.scala 151:92:@13375.4]
  wire  _T_15417; // @[LoadQueue.scala 152:41:@13376.4]
  wire  _T_15418; // @[LoadQueue.scala 153:30:@13377.4]
  wire  conflict_13_8; // @[LoadQueue.scala 152:68:@13378.4]
  wire  _T_15420; // @[LoadQueue.scala 151:92:@13380.4]
  wire  _T_15421; // @[LoadQueue.scala 152:41:@13381.4]
  wire  _T_15422; // @[LoadQueue.scala 153:30:@13382.4]
  wire  conflict_13_9; // @[LoadQueue.scala 152:68:@13383.4]
  wire  _T_15424; // @[LoadQueue.scala 151:92:@13385.4]
  wire  _T_15425; // @[LoadQueue.scala 152:41:@13386.4]
  wire  _T_15426; // @[LoadQueue.scala 153:30:@13387.4]
  wire  conflict_13_10; // @[LoadQueue.scala 152:68:@13388.4]
  wire  _T_15428; // @[LoadQueue.scala 151:92:@13390.4]
  wire  _T_15429; // @[LoadQueue.scala 152:41:@13391.4]
  wire  _T_15430; // @[LoadQueue.scala 153:30:@13392.4]
  wire  conflict_13_11; // @[LoadQueue.scala 152:68:@13393.4]
  wire  _T_15432; // @[LoadQueue.scala 151:92:@13395.4]
  wire  _T_15433; // @[LoadQueue.scala 152:41:@13396.4]
  wire  _T_15434; // @[LoadQueue.scala 153:30:@13397.4]
  wire  conflict_13_12; // @[LoadQueue.scala 152:68:@13398.4]
  wire  _T_15436; // @[LoadQueue.scala 151:92:@13400.4]
  wire  _T_15437; // @[LoadQueue.scala 152:41:@13401.4]
  wire  _T_15438; // @[LoadQueue.scala 153:30:@13402.4]
  wire  conflict_13_13; // @[LoadQueue.scala 152:68:@13403.4]
  wire  _T_15440; // @[LoadQueue.scala 151:92:@13405.4]
  wire  _T_15441; // @[LoadQueue.scala 152:41:@13406.4]
  wire  _T_15442; // @[LoadQueue.scala 153:30:@13407.4]
  wire  conflict_13_14; // @[LoadQueue.scala 152:68:@13408.4]
  wire  _T_15444; // @[LoadQueue.scala 151:92:@13410.4]
  wire  _T_15445; // @[LoadQueue.scala 152:41:@13411.4]
  wire  _T_15446; // @[LoadQueue.scala 153:30:@13412.4]
  wire  conflict_13_15; // @[LoadQueue.scala 152:68:@13413.4]
  wire  _T_15448; // @[LoadQueue.scala 151:92:@13415.4]
  wire  _T_15449; // @[LoadQueue.scala 152:41:@13416.4]
  wire  _T_15450; // @[LoadQueue.scala 153:30:@13417.4]
  wire  conflict_14_0; // @[LoadQueue.scala 152:68:@13418.4]
  wire  _T_15452; // @[LoadQueue.scala 151:92:@13420.4]
  wire  _T_15453; // @[LoadQueue.scala 152:41:@13421.4]
  wire  _T_15454; // @[LoadQueue.scala 153:30:@13422.4]
  wire  conflict_14_1; // @[LoadQueue.scala 152:68:@13423.4]
  wire  _T_15456; // @[LoadQueue.scala 151:92:@13425.4]
  wire  _T_15457; // @[LoadQueue.scala 152:41:@13426.4]
  wire  _T_15458; // @[LoadQueue.scala 153:30:@13427.4]
  wire  conflict_14_2; // @[LoadQueue.scala 152:68:@13428.4]
  wire  _T_15460; // @[LoadQueue.scala 151:92:@13430.4]
  wire  _T_15461; // @[LoadQueue.scala 152:41:@13431.4]
  wire  _T_15462; // @[LoadQueue.scala 153:30:@13432.4]
  wire  conflict_14_3; // @[LoadQueue.scala 152:68:@13433.4]
  wire  _T_15464; // @[LoadQueue.scala 151:92:@13435.4]
  wire  _T_15465; // @[LoadQueue.scala 152:41:@13436.4]
  wire  _T_15466; // @[LoadQueue.scala 153:30:@13437.4]
  wire  conflict_14_4; // @[LoadQueue.scala 152:68:@13438.4]
  wire  _T_15468; // @[LoadQueue.scala 151:92:@13440.4]
  wire  _T_15469; // @[LoadQueue.scala 152:41:@13441.4]
  wire  _T_15470; // @[LoadQueue.scala 153:30:@13442.4]
  wire  conflict_14_5; // @[LoadQueue.scala 152:68:@13443.4]
  wire  _T_15472; // @[LoadQueue.scala 151:92:@13445.4]
  wire  _T_15473; // @[LoadQueue.scala 152:41:@13446.4]
  wire  _T_15474; // @[LoadQueue.scala 153:30:@13447.4]
  wire  conflict_14_6; // @[LoadQueue.scala 152:68:@13448.4]
  wire  _T_15476; // @[LoadQueue.scala 151:92:@13450.4]
  wire  _T_15477; // @[LoadQueue.scala 152:41:@13451.4]
  wire  _T_15478; // @[LoadQueue.scala 153:30:@13452.4]
  wire  conflict_14_7; // @[LoadQueue.scala 152:68:@13453.4]
  wire  _T_15480; // @[LoadQueue.scala 151:92:@13455.4]
  wire  _T_15481; // @[LoadQueue.scala 152:41:@13456.4]
  wire  _T_15482; // @[LoadQueue.scala 153:30:@13457.4]
  wire  conflict_14_8; // @[LoadQueue.scala 152:68:@13458.4]
  wire  _T_15484; // @[LoadQueue.scala 151:92:@13460.4]
  wire  _T_15485; // @[LoadQueue.scala 152:41:@13461.4]
  wire  _T_15486; // @[LoadQueue.scala 153:30:@13462.4]
  wire  conflict_14_9; // @[LoadQueue.scala 152:68:@13463.4]
  wire  _T_15488; // @[LoadQueue.scala 151:92:@13465.4]
  wire  _T_15489; // @[LoadQueue.scala 152:41:@13466.4]
  wire  _T_15490; // @[LoadQueue.scala 153:30:@13467.4]
  wire  conflict_14_10; // @[LoadQueue.scala 152:68:@13468.4]
  wire  _T_15492; // @[LoadQueue.scala 151:92:@13470.4]
  wire  _T_15493; // @[LoadQueue.scala 152:41:@13471.4]
  wire  _T_15494; // @[LoadQueue.scala 153:30:@13472.4]
  wire  conflict_14_11; // @[LoadQueue.scala 152:68:@13473.4]
  wire  _T_15496; // @[LoadQueue.scala 151:92:@13475.4]
  wire  _T_15497; // @[LoadQueue.scala 152:41:@13476.4]
  wire  _T_15498; // @[LoadQueue.scala 153:30:@13477.4]
  wire  conflict_14_12; // @[LoadQueue.scala 152:68:@13478.4]
  wire  _T_15500; // @[LoadQueue.scala 151:92:@13480.4]
  wire  _T_15501; // @[LoadQueue.scala 152:41:@13481.4]
  wire  _T_15502; // @[LoadQueue.scala 153:30:@13482.4]
  wire  conflict_14_13; // @[LoadQueue.scala 152:68:@13483.4]
  wire  _T_15504; // @[LoadQueue.scala 151:92:@13485.4]
  wire  _T_15505; // @[LoadQueue.scala 152:41:@13486.4]
  wire  _T_15506; // @[LoadQueue.scala 153:30:@13487.4]
  wire  conflict_14_14; // @[LoadQueue.scala 152:68:@13488.4]
  wire  _T_15508; // @[LoadQueue.scala 151:92:@13490.4]
  wire  _T_15509; // @[LoadQueue.scala 152:41:@13491.4]
  wire  _T_15510; // @[LoadQueue.scala 153:30:@13492.4]
  wire  conflict_14_15; // @[LoadQueue.scala 152:68:@13493.4]
  wire  _T_15512; // @[LoadQueue.scala 151:92:@13495.4]
  wire  _T_15513; // @[LoadQueue.scala 152:41:@13496.4]
  wire  _T_15514; // @[LoadQueue.scala 153:30:@13497.4]
  wire  conflict_15_0; // @[LoadQueue.scala 152:68:@13498.4]
  wire  _T_15516; // @[LoadQueue.scala 151:92:@13500.4]
  wire  _T_15517; // @[LoadQueue.scala 152:41:@13501.4]
  wire  _T_15518; // @[LoadQueue.scala 153:30:@13502.4]
  wire  conflict_15_1; // @[LoadQueue.scala 152:68:@13503.4]
  wire  _T_15520; // @[LoadQueue.scala 151:92:@13505.4]
  wire  _T_15521; // @[LoadQueue.scala 152:41:@13506.4]
  wire  _T_15522; // @[LoadQueue.scala 153:30:@13507.4]
  wire  conflict_15_2; // @[LoadQueue.scala 152:68:@13508.4]
  wire  _T_15524; // @[LoadQueue.scala 151:92:@13510.4]
  wire  _T_15525; // @[LoadQueue.scala 152:41:@13511.4]
  wire  _T_15526; // @[LoadQueue.scala 153:30:@13512.4]
  wire  conflict_15_3; // @[LoadQueue.scala 152:68:@13513.4]
  wire  _T_15528; // @[LoadQueue.scala 151:92:@13515.4]
  wire  _T_15529; // @[LoadQueue.scala 152:41:@13516.4]
  wire  _T_15530; // @[LoadQueue.scala 153:30:@13517.4]
  wire  conflict_15_4; // @[LoadQueue.scala 152:68:@13518.4]
  wire  _T_15532; // @[LoadQueue.scala 151:92:@13520.4]
  wire  _T_15533; // @[LoadQueue.scala 152:41:@13521.4]
  wire  _T_15534; // @[LoadQueue.scala 153:30:@13522.4]
  wire  conflict_15_5; // @[LoadQueue.scala 152:68:@13523.4]
  wire  _T_15536; // @[LoadQueue.scala 151:92:@13525.4]
  wire  _T_15537; // @[LoadQueue.scala 152:41:@13526.4]
  wire  _T_15538; // @[LoadQueue.scala 153:30:@13527.4]
  wire  conflict_15_6; // @[LoadQueue.scala 152:68:@13528.4]
  wire  _T_15540; // @[LoadQueue.scala 151:92:@13530.4]
  wire  _T_15541; // @[LoadQueue.scala 152:41:@13531.4]
  wire  _T_15542; // @[LoadQueue.scala 153:30:@13532.4]
  wire  conflict_15_7; // @[LoadQueue.scala 152:68:@13533.4]
  wire  _T_15544; // @[LoadQueue.scala 151:92:@13535.4]
  wire  _T_15545; // @[LoadQueue.scala 152:41:@13536.4]
  wire  _T_15546; // @[LoadQueue.scala 153:30:@13537.4]
  wire  conflict_15_8; // @[LoadQueue.scala 152:68:@13538.4]
  wire  _T_15548; // @[LoadQueue.scala 151:92:@13540.4]
  wire  _T_15549; // @[LoadQueue.scala 152:41:@13541.4]
  wire  _T_15550; // @[LoadQueue.scala 153:30:@13542.4]
  wire  conflict_15_9; // @[LoadQueue.scala 152:68:@13543.4]
  wire  _T_15552; // @[LoadQueue.scala 151:92:@13545.4]
  wire  _T_15553; // @[LoadQueue.scala 152:41:@13546.4]
  wire  _T_15554; // @[LoadQueue.scala 153:30:@13547.4]
  wire  conflict_15_10; // @[LoadQueue.scala 152:68:@13548.4]
  wire  _T_15556; // @[LoadQueue.scala 151:92:@13550.4]
  wire  _T_15557; // @[LoadQueue.scala 152:41:@13551.4]
  wire  _T_15558; // @[LoadQueue.scala 153:30:@13552.4]
  wire  conflict_15_11; // @[LoadQueue.scala 152:68:@13553.4]
  wire  _T_15560; // @[LoadQueue.scala 151:92:@13555.4]
  wire  _T_15561; // @[LoadQueue.scala 152:41:@13556.4]
  wire  _T_15562; // @[LoadQueue.scala 153:30:@13557.4]
  wire  conflict_15_12; // @[LoadQueue.scala 152:68:@13558.4]
  wire  _T_15564; // @[LoadQueue.scala 151:92:@13560.4]
  wire  _T_15565; // @[LoadQueue.scala 152:41:@13561.4]
  wire  _T_15566; // @[LoadQueue.scala 153:30:@13562.4]
  wire  conflict_15_13; // @[LoadQueue.scala 152:68:@13563.4]
  wire  _T_15568; // @[LoadQueue.scala 151:92:@13565.4]
  wire  _T_15569; // @[LoadQueue.scala 152:41:@13566.4]
  wire  _T_15570; // @[LoadQueue.scala 153:30:@13567.4]
  wire  conflict_15_14; // @[LoadQueue.scala 152:68:@13568.4]
  wire  _T_15572; // @[LoadQueue.scala 151:92:@13570.4]
  wire  _T_15573; // @[LoadQueue.scala 152:41:@13571.4]
  wire  _T_15574; // @[LoadQueue.scala 153:30:@13572.4]
  wire  conflict_15_15; // @[LoadQueue.scala 152:68:@13573.4]
  wire  _T_16807; // @[LoadQueue.scala 163:13:@13576.4]
  wire  storeAddrNotKnownFlags_0_0; // @[LoadQueue.scala 163:19:@13577.4]
  wire  _T_16810; // @[LoadQueue.scala 163:13:@13578.4]
  wire  storeAddrNotKnownFlags_0_1; // @[LoadQueue.scala 163:19:@13579.4]
  wire  _T_16813; // @[LoadQueue.scala 163:13:@13580.4]
  wire  storeAddrNotKnownFlags_0_2; // @[LoadQueue.scala 163:19:@13581.4]
  wire  _T_16816; // @[LoadQueue.scala 163:13:@13582.4]
  wire  storeAddrNotKnownFlags_0_3; // @[LoadQueue.scala 163:19:@13583.4]
  wire  _T_16819; // @[LoadQueue.scala 163:13:@13584.4]
  wire  storeAddrNotKnownFlags_0_4; // @[LoadQueue.scala 163:19:@13585.4]
  wire  _T_16822; // @[LoadQueue.scala 163:13:@13586.4]
  wire  storeAddrNotKnownFlags_0_5; // @[LoadQueue.scala 163:19:@13587.4]
  wire  _T_16825; // @[LoadQueue.scala 163:13:@13588.4]
  wire  storeAddrNotKnownFlags_0_6; // @[LoadQueue.scala 163:19:@13589.4]
  wire  _T_16828; // @[LoadQueue.scala 163:13:@13590.4]
  wire  storeAddrNotKnownFlags_0_7; // @[LoadQueue.scala 163:19:@13591.4]
  wire  _T_16831; // @[LoadQueue.scala 163:13:@13592.4]
  wire  storeAddrNotKnownFlags_0_8; // @[LoadQueue.scala 163:19:@13593.4]
  wire  _T_16834; // @[LoadQueue.scala 163:13:@13594.4]
  wire  storeAddrNotKnownFlags_0_9; // @[LoadQueue.scala 163:19:@13595.4]
  wire  _T_16837; // @[LoadQueue.scala 163:13:@13596.4]
  wire  storeAddrNotKnownFlags_0_10; // @[LoadQueue.scala 163:19:@13597.4]
  wire  _T_16840; // @[LoadQueue.scala 163:13:@13598.4]
  wire  storeAddrNotKnownFlags_0_11; // @[LoadQueue.scala 163:19:@13599.4]
  wire  _T_16843; // @[LoadQueue.scala 163:13:@13600.4]
  wire  storeAddrNotKnownFlags_0_12; // @[LoadQueue.scala 163:19:@13601.4]
  wire  _T_16846; // @[LoadQueue.scala 163:13:@13602.4]
  wire  storeAddrNotKnownFlags_0_13; // @[LoadQueue.scala 163:19:@13603.4]
  wire  _T_16849; // @[LoadQueue.scala 163:13:@13604.4]
  wire  storeAddrNotKnownFlags_0_14; // @[LoadQueue.scala 163:19:@13605.4]
  wire  _T_16852; // @[LoadQueue.scala 163:13:@13606.4]
  wire  storeAddrNotKnownFlags_0_15; // @[LoadQueue.scala 163:19:@13607.4]
  wire  storeAddrNotKnownFlags_1_0; // @[LoadQueue.scala 163:19:@13625.4]
  wire  storeAddrNotKnownFlags_1_1; // @[LoadQueue.scala 163:19:@13627.4]
  wire  storeAddrNotKnownFlags_1_2; // @[LoadQueue.scala 163:19:@13629.4]
  wire  storeAddrNotKnownFlags_1_3; // @[LoadQueue.scala 163:19:@13631.4]
  wire  storeAddrNotKnownFlags_1_4; // @[LoadQueue.scala 163:19:@13633.4]
  wire  storeAddrNotKnownFlags_1_5; // @[LoadQueue.scala 163:19:@13635.4]
  wire  storeAddrNotKnownFlags_1_6; // @[LoadQueue.scala 163:19:@13637.4]
  wire  storeAddrNotKnownFlags_1_7; // @[LoadQueue.scala 163:19:@13639.4]
  wire  storeAddrNotKnownFlags_1_8; // @[LoadQueue.scala 163:19:@13641.4]
  wire  storeAddrNotKnownFlags_1_9; // @[LoadQueue.scala 163:19:@13643.4]
  wire  storeAddrNotKnownFlags_1_10; // @[LoadQueue.scala 163:19:@13645.4]
  wire  storeAddrNotKnownFlags_1_11; // @[LoadQueue.scala 163:19:@13647.4]
  wire  storeAddrNotKnownFlags_1_12; // @[LoadQueue.scala 163:19:@13649.4]
  wire  storeAddrNotKnownFlags_1_13; // @[LoadQueue.scala 163:19:@13651.4]
  wire  storeAddrNotKnownFlags_1_14; // @[LoadQueue.scala 163:19:@13653.4]
  wire  storeAddrNotKnownFlags_1_15; // @[LoadQueue.scala 163:19:@13655.4]
  wire  storeAddrNotKnownFlags_2_0; // @[LoadQueue.scala 163:19:@13673.4]
  wire  storeAddrNotKnownFlags_2_1; // @[LoadQueue.scala 163:19:@13675.4]
  wire  storeAddrNotKnownFlags_2_2; // @[LoadQueue.scala 163:19:@13677.4]
  wire  storeAddrNotKnownFlags_2_3; // @[LoadQueue.scala 163:19:@13679.4]
  wire  storeAddrNotKnownFlags_2_4; // @[LoadQueue.scala 163:19:@13681.4]
  wire  storeAddrNotKnownFlags_2_5; // @[LoadQueue.scala 163:19:@13683.4]
  wire  storeAddrNotKnownFlags_2_6; // @[LoadQueue.scala 163:19:@13685.4]
  wire  storeAddrNotKnownFlags_2_7; // @[LoadQueue.scala 163:19:@13687.4]
  wire  storeAddrNotKnownFlags_2_8; // @[LoadQueue.scala 163:19:@13689.4]
  wire  storeAddrNotKnownFlags_2_9; // @[LoadQueue.scala 163:19:@13691.4]
  wire  storeAddrNotKnownFlags_2_10; // @[LoadQueue.scala 163:19:@13693.4]
  wire  storeAddrNotKnownFlags_2_11; // @[LoadQueue.scala 163:19:@13695.4]
  wire  storeAddrNotKnownFlags_2_12; // @[LoadQueue.scala 163:19:@13697.4]
  wire  storeAddrNotKnownFlags_2_13; // @[LoadQueue.scala 163:19:@13699.4]
  wire  storeAddrNotKnownFlags_2_14; // @[LoadQueue.scala 163:19:@13701.4]
  wire  storeAddrNotKnownFlags_2_15; // @[LoadQueue.scala 163:19:@13703.4]
  wire  storeAddrNotKnownFlags_3_0; // @[LoadQueue.scala 163:19:@13721.4]
  wire  storeAddrNotKnownFlags_3_1; // @[LoadQueue.scala 163:19:@13723.4]
  wire  storeAddrNotKnownFlags_3_2; // @[LoadQueue.scala 163:19:@13725.4]
  wire  storeAddrNotKnownFlags_3_3; // @[LoadQueue.scala 163:19:@13727.4]
  wire  storeAddrNotKnownFlags_3_4; // @[LoadQueue.scala 163:19:@13729.4]
  wire  storeAddrNotKnownFlags_3_5; // @[LoadQueue.scala 163:19:@13731.4]
  wire  storeAddrNotKnownFlags_3_6; // @[LoadQueue.scala 163:19:@13733.4]
  wire  storeAddrNotKnownFlags_3_7; // @[LoadQueue.scala 163:19:@13735.4]
  wire  storeAddrNotKnownFlags_3_8; // @[LoadQueue.scala 163:19:@13737.4]
  wire  storeAddrNotKnownFlags_3_9; // @[LoadQueue.scala 163:19:@13739.4]
  wire  storeAddrNotKnownFlags_3_10; // @[LoadQueue.scala 163:19:@13741.4]
  wire  storeAddrNotKnownFlags_3_11; // @[LoadQueue.scala 163:19:@13743.4]
  wire  storeAddrNotKnownFlags_3_12; // @[LoadQueue.scala 163:19:@13745.4]
  wire  storeAddrNotKnownFlags_3_13; // @[LoadQueue.scala 163:19:@13747.4]
  wire  storeAddrNotKnownFlags_3_14; // @[LoadQueue.scala 163:19:@13749.4]
  wire  storeAddrNotKnownFlags_3_15; // @[LoadQueue.scala 163:19:@13751.4]
  wire  storeAddrNotKnownFlags_4_0; // @[LoadQueue.scala 163:19:@13769.4]
  wire  storeAddrNotKnownFlags_4_1; // @[LoadQueue.scala 163:19:@13771.4]
  wire  storeAddrNotKnownFlags_4_2; // @[LoadQueue.scala 163:19:@13773.4]
  wire  storeAddrNotKnownFlags_4_3; // @[LoadQueue.scala 163:19:@13775.4]
  wire  storeAddrNotKnownFlags_4_4; // @[LoadQueue.scala 163:19:@13777.4]
  wire  storeAddrNotKnownFlags_4_5; // @[LoadQueue.scala 163:19:@13779.4]
  wire  storeAddrNotKnownFlags_4_6; // @[LoadQueue.scala 163:19:@13781.4]
  wire  storeAddrNotKnownFlags_4_7; // @[LoadQueue.scala 163:19:@13783.4]
  wire  storeAddrNotKnownFlags_4_8; // @[LoadQueue.scala 163:19:@13785.4]
  wire  storeAddrNotKnownFlags_4_9; // @[LoadQueue.scala 163:19:@13787.4]
  wire  storeAddrNotKnownFlags_4_10; // @[LoadQueue.scala 163:19:@13789.4]
  wire  storeAddrNotKnownFlags_4_11; // @[LoadQueue.scala 163:19:@13791.4]
  wire  storeAddrNotKnownFlags_4_12; // @[LoadQueue.scala 163:19:@13793.4]
  wire  storeAddrNotKnownFlags_4_13; // @[LoadQueue.scala 163:19:@13795.4]
  wire  storeAddrNotKnownFlags_4_14; // @[LoadQueue.scala 163:19:@13797.4]
  wire  storeAddrNotKnownFlags_4_15; // @[LoadQueue.scala 163:19:@13799.4]
  wire  storeAddrNotKnownFlags_5_0; // @[LoadQueue.scala 163:19:@13817.4]
  wire  storeAddrNotKnownFlags_5_1; // @[LoadQueue.scala 163:19:@13819.4]
  wire  storeAddrNotKnownFlags_5_2; // @[LoadQueue.scala 163:19:@13821.4]
  wire  storeAddrNotKnownFlags_5_3; // @[LoadQueue.scala 163:19:@13823.4]
  wire  storeAddrNotKnownFlags_5_4; // @[LoadQueue.scala 163:19:@13825.4]
  wire  storeAddrNotKnownFlags_5_5; // @[LoadQueue.scala 163:19:@13827.4]
  wire  storeAddrNotKnownFlags_5_6; // @[LoadQueue.scala 163:19:@13829.4]
  wire  storeAddrNotKnownFlags_5_7; // @[LoadQueue.scala 163:19:@13831.4]
  wire  storeAddrNotKnownFlags_5_8; // @[LoadQueue.scala 163:19:@13833.4]
  wire  storeAddrNotKnownFlags_5_9; // @[LoadQueue.scala 163:19:@13835.4]
  wire  storeAddrNotKnownFlags_5_10; // @[LoadQueue.scala 163:19:@13837.4]
  wire  storeAddrNotKnownFlags_5_11; // @[LoadQueue.scala 163:19:@13839.4]
  wire  storeAddrNotKnownFlags_5_12; // @[LoadQueue.scala 163:19:@13841.4]
  wire  storeAddrNotKnownFlags_5_13; // @[LoadQueue.scala 163:19:@13843.4]
  wire  storeAddrNotKnownFlags_5_14; // @[LoadQueue.scala 163:19:@13845.4]
  wire  storeAddrNotKnownFlags_5_15; // @[LoadQueue.scala 163:19:@13847.4]
  wire  storeAddrNotKnownFlags_6_0; // @[LoadQueue.scala 163:19:@13865.4]
  wire  storeAddrNotKnownFlags_6_1; // @[LoadQueue.scala 163:19:@13867.4]
  wire  storeAddrNotKnownFlags_6_2; // @[LoadQueue.scala 163:19:@13869.4]
  wire  storeAddrNotKnownFlags_6_3; // @[LoadQueue.scala 163:19:@13871.4]
  wire  storeAddrNotKnownFlags_6_4; // @[LoadQueue.scala 163:19:@13873.4]
  wire  storeAddrNotKnownFlags_6_5; // @[LoadQueue.scala 163:19:@13875.4]
  wire  storeAddrNotKnownFlags_6_6; // @[LoadQueue.scala 163:19:@13877.4]
  wire  storeAddrNotKnownFlags_6_7; // @[LoadQueue.scala 163:19:@13879.4]
  wire  storeAddrNotKnownFlags_6_8; // @[LoadQueue.scala 163:19:@13881.4]
  wire  storeAddrNotKnownFlags_6_9; // @[LoadQueue.scala 163:19:@13883.4]
  wire  storeAddrNotKnownFlags_6_10; // @[LoadQueue.scala 163:19:@13885.4]
  wire  storeAddrNotKnownFlags_6_11; // @[LoadQueue.scala 163:19:@13887.4]
  wire  storeAddrNotKnownFlags_6_12; // @[LoadQueue.scala 163:19:@13889.4]
  wire  storeAddrNotKnownFlags_6_13; // @[LoadQueue.scala 163:19:@13891.4]
  wire  storeAddrNotKnownFlags_6_14; // @[LoadQueue.scala 163:19:@13893.4]
  wire  storeAddrNotKnownFlags_6_15; // @[LoadQueue.scala 163:19:@13895.4]
  wire  storeAddrNotKnownFlags_7_0; // @[LoadQueue.scala 163:19:@13913.4]
  wire  storeAddrNotKnownFlags_7_1; // @[LoadQueue.scala 163:19:@13915.4]
  wire  storeAddrNotKnownFlags_7_2; // @[LoadQueue.scala 163:19:@13917.4]
  wire  storeAddrNotKnownFlags_7_3; // @[LoadQueue.scala 163:19:@13919.4]
  wire  storeAddrNotKnownFlags_7_4; // @[LoadQueue.scala 163:19:@13921.4]
  wire  storeAddrNotKnownFlags_7_5; // @[LoadQueue.scala 163:19:@13923.4]
  wire  storeAddrNotKnownFlags_7_6; // @[LoadQueue.scala 163:19:@13925.4]
  wire  storeAddrNotKnownFlags_7_7; // @[LoadQueue.scala 163:19:@13927.4]
  wire  storeAddrNotKnownFlags_7_8; // @[LoadQueue.scala 163:19:@13929.4]
  wire  storeAddrNotKnownFlags_7_9; // @[LoadQueue.scala 163:19:@13931.4]
  wire  storeAddrNotKnownFlags_7_10; // @[LoadQueue.scala 163:19:@13933.4]
  wire  storeAddrNotKnownFlags_7_11; // @[LoadQueue.scala 163:19:@13935.4]
  wire  storeAddrNotKnownFlags_7_12; // @[LoadQueue.scala 163:19:@13937.4]
  wire  storeAddrNotKnownFlags_7_13; // @[LoadQueue.scala 163:19:@13939.4]
  wire  storeAddrNotKnownFlags_7_14; // @[LoadQueue.scala 163:19:@13941.4]
  wire  storeAddrNotKnownFlags_7_15; // @[LoadQueue.scala 163:19:@13943.4]
  wire  storeAddrNotKnownFlags_8_0; // @[LoadQueue.scala 163:19:@13961.4]
  wire  storeAddrNotKnownFlags_8_1; // @[LoadQueue.scala 163:19:@13963.4]
  wire  storeAddrNotKnownFlags_8_2; // @[LoadQueue.scala 163:19:@13965.4]
  wire  storeAddrNotKnownFlags_8_3; // @[LoadQueue.scala 163:19:@13967.4]
  wire  storeAddrNotKnownFlags_8_4; // @[LoadQueue.scala 163:19:@13969.4]
  wire  storeAddrNotKnownFlags_8_5; // @[LoadQueue.scala 163:19:@13971.4]
  wire  storeAddrNotKnownFlags_8_6; // @[LoadQueue.scala 163:19:@13973.4]
  wire  storeAddrNotKnownFlags_8_7; // @[LoadQueue.scala 163:19:@13975.4]
  wire  storeAddrNotKnownFlags_8_8; // @[LoadQueue.scala 163:19:@13977.4]
  wire  storeAddrNotKnownFlags_8_9; // @[LoadQueue.scala 163:19:@13979.4]
  wire  storeAddrNotKnownFlags_8_10; // @[LoadQueue.scala 163:19:@13981.4]
  wire  storeAddrNotKnownFlags_8_11; // @[LoadQueue.scala 163:19:@13983.4]
  wire  storeAddrNotKnownFlags_8_12; // @[LoadQueue.scala 163:19:@13985.4]
  wire  storeAddrNotKnownFlags_8_13; // @[LoadQueue.scala 163:19:@13987.4]
  wire  storeAddrNotKnownFlags_8_14; // @[LoadQueue.scala 163:19:@13989.4]
  wire  storeAddrNotKnownFlags_8_15; // @[LoadQueue.scala 163:19:@13991.4]
  wire  storeAddrNotKnownFlags_9_0; // @[LoadQueue.scala 163:19:@14009.4]
  wire  storeAddrNotKnownFlags_9_1; // @[LoadQueue.scala 163:19:@14011.4]
  wire  storeAddrNotKnownFlags_9_2; // @[LoadQueue.scala 163:19:@14013.4]
  wire  storeAddrNotKnownFlags_9_3; // @[LoadQueue.scala 163:19:@14015.4]
  wire  storeAddrNotKnownFlags_9_4; // @[LoadQueue.scala 163:19:@14017.4]
  wire  storeAddrNotKnownFlags_9_5; // @[LoadQueue.scala 163:19:@14019.4]
  wire  storeAddrNotKnownFlags_9_6; // @[LoadQueue.scala 163:19:@14021.4]
  wire  storeAddrNotKnownFlags_9_7; // @[LoadQueue.scala 163:19:@14023.4]
  wire  storeAddrNotKnownFlags_9_8; // @[LoadQueue.scala 163:19:@14025.4]
  wire  storeAddrNotKnownFlags_9_9; // @[LoadQueue.scala 163:19:@14027.4]
  wire  storeAddrNotKnownFlags_9_10; // @[LoadQueue.scala 163:19:@14029.4]
  wire  storeAddrNotKnownFlags_9_11; // @[LoadQueue.scala 163:19:@14031.4]
  wire  storeAddrNotKnownFlags_9_12; // @[LoadQueue.scala 163:19:@14033.4]
  wire  storeAddrNotKnownFlags_9_13; // @[LoadQueue.scala 163:19:@14035.4]
  wire  storeAddrNotKnownFlags_9_14; // @[LoadQueue.scala 163:19:@14037.4]
  wire  storeAddrNotKnownFlags_9_15; // @[LoadQueue.scala 163:19:@14039.4]
  wire  storeAddrNotKnownFlags_10_0; // @[LoadQueue.scala 163:19:@14057.4]
  wire  storeAddrNotKnownFlags_10_1; // @[LoadQueue.scala 163:19:@14059.4]
  wire  storeAddrNotKnownFlags_10_2; // @[LoadQueue.scala 163:19:@14061.4]
  wire  storeAddrNotKnownFlags_10_3; // @[LoadQueue.scala 163:19:@14063.4]
  wire  storeAddrNotKnownFlags_10_4; // @[LoadQueue.scala 163:19:@14065.4]
  wire  storeAddrNotKnownFlags_10_5; // @[LoadQueue.scala 163:19:@14067.4]
  wire  storeAddrNotKnownFlags_10_6; // @[LoadQueue.scala 163:19:@14069.4]
  wire  storeAddrNotKnownFlags_10_7; // @[LoadQueue.scala 163:19:@14071.4]
  wire  storeAddrNotKnownFlags_10_8; // @[LoadQueue.scala 163:19:@14073.4]
  wire  storeAddrNotKnownFlags_10_9; // @[LoadQueue.scala 163:19:@14075.4]
  wire  storeAddrNotKnownFlags_10_10; // @[LoadQueue.scala 163:19:@14077.4]
  wire  storeAddrNotKnownFlags_10_11; // @[LoadQueue.scala 163:19:@14079.4]
  wire  storeAddrNotKnownFlags_10_12; // @[LoadQueue.scala 163:19:@14081.4]
  wire  storeAddrNotKnownFlags_10_13; // @[LoadQueue.scala 163:19:@14083.4]
  wire  storeAddrNotKnownFlags_10_14; // @[LoadQueue.scala 163:19:@14085.4]
  wire  storeAddrNotKnownFlags_10_15; // @[LoadQueue.scala 163:19:@14087.4]
  wire  storeAddrNotKnownFlags_11_0; // @[LoadQueue.scala 163:19:@14105.4]
  wire  storeAddrNotKnownFlags_11_1; // @[LoadQueue.scala 163:19:@14107.4]
  wire  storeAddrNotKnownFlags_11_2; // @[LoadQueue.scala 163:19:@14109.4]
  wire  storeAddrNotKnownFlags_11_3; // @[LoadQueue.scala 163:19:@14111.4]
  wire  storeAddrNotKnownFlags_11_4; // @[LoadQueue.scala 163:19:@14113.4]
  wire  storeAddrNotKnownFlags_11_5; // @[LoadQueue.scala 163:19:@14115.4]
  wire  storeAddrNotKnownFlags_11_6; // @[LoadQueue.scala 163:19:@14117.4]
  wire  storeAddrNotKnownFlags_11_7; // @[LoadQueue.scala 163:19:@14119.4]
  wire  storeAddrNotKnownFlags_11_8; // @[LoadQueue.scala 163:19:@14121.4]
  wire  storeAddrNotKnownFlags_11_9; // @[LoadQueue.scala 163:19:@14123.4]
  wire  storeAddrNotKnownFlags_11_10; // @[LoadQueue.scala 163:19:@14125.4]
  wire  storeAddrNotKnownFlags_11_11; // @[LoadQueue.scala 163:19:@14127.4]
  wire  storeAddrNotKnownFlags_11_12; // @[LoadQueue.scala 163:19:@14129.4]
  wire  storeAddrNotKnownFlags_11_13; // @[LoadQueue.scala 163:19:@14131.4]
  wire  storeAddrNotKnownFlags_11_14; // @[LoadQueue.scala 163:19:@14133.4]
  wire  storeAddrNotKnownFlags_11_15; // @[LoadQueue.scala 163:19:@14135.4]
  wire  storeAddrNotKnownFlags_12_0; // @[LoadQueue.scala 163:19:@14153.4]
  wire  storeAddrNotKnownFlags_12_1; // @[LoadQueue.scala 163:19:@14155.4]
  wire  storeAddrNotKnownFlags_12_2; // @[LoadQueue.scala 163:19:@14157.4]
  wire  storeAddrNotKnownFlags_12_3; // @[LoadQueue.scala 163:19:@14159.4]
  wire  storeAddrNotKnownFlags_12_4; // @[LoadQueue.scala 163:19:@14161.4]
  wire  storeAddrNotKnownFlags_12_5; // @[LoadQueue.scala 163:19:@14163.4]
  wire  storeAddrNotKnownFlags_12_6; // @[LoadQueue.scala 163:19:@14165.4]
  wire  storeAddrNotKnownFlags_12_7; // @[LoadQueue.scala 163:19:@14167.4]
  wire  storeAddrNotKnownFlags_12_8; // @[LoadQueue.scala 163:19:@14169.4]
  wire  storeAddrNotKnownFlags_12_9; // @[LoadQueue.scala 163:19:@14171.4]
  wire  storeAddrNotKnownFlags_12_10; // @[LoadQueue.scala 163:19:@14173.4]
  wire  storeAddrNotKnownFlags_12_11; // @[LoadQueue.scala 163:19:@14175.4]
  wire  storeAddrNotKnownFlags_12_12; // @[LoadQueue.scala 163:19:@14177.4]
  wire  storeAddrNotKnownFlags_12_13; // @[LoadQueue.scala 163:19:@14179.4]
  wire  storeAddrNotKnownFlags_12_14; // @[LoadQueue.scala 163:19:@14181.4]
  wire  storeAddrNotKnownFlags_12_15; // @[LoadQueue.scala 163:19:@14183.4]
  wire  storeAddrNotKnownFlags_13_0; // @[LoadQueue.scala 163:19:@14201.4]
  wire  storeAddrNotKnownFlags_13_1; // @[LoadQueue.scala 163:19:@14203.4]
  wire  storeAddrNotKnownFlags_13_2; // @[LoadQueue.scala 163:19:@14205.4]
  wire  storeAddrNotKnownFlags_13_3; // @[LoadQueue.scala 163:19:@14207.4]
  wire  storeAddrNotKnownFlags_13_4; // @[LoadQueue.scala 163:19:@14209.4]
  wire  storeAddrNotKnownFlags_13_5; // @[LoadQueue.scala 163:19:@14211.4]
  wire  storeAddrNotKnownFlags_13_6; // @[LoadQueue.scala 163:19:@14213.4]
  wire  storeAddrNotKnownFlags_13_7; // @[LoadQueue.scala 163:19:@14215.4]
  wire  storeAddrNotKnownFlags_13_8; // @[LoadQueue.scala 163:19:@14217.4]
  wire  storeAddrNotKnownFlags_13_9; // @[LoadQueue.scala 163:19:@14219.4]
  wire  storeAddrNotKnownFlags_13_10; // @[LoadQueue.scala 163:19:@14221.4]
  wire  storeAddrNotKnownFlags_13_11; // @[LoadQueue.scala 163:19:@14223.4]
  wire  storeAddrNotKnownFlags_13_12; // @[LoadQueue.scala 163:19:@14225.4]
  wire  storeAddrNotKnownFlags_13_13; // @[LoadQueue.scala 163:19:@14227.4]
  wire  storeAddrNotKnownFlags_13_14; // @[LoadQueue.scala 163:19:@14229.4]
  wire  storeAddrNotKnownFlags_13_15; // @[LoadQueue.scala 163:19:@14231.4]
  wire  storeAddrNotKnownFlags_14_0; // @[LoadQueue.scala 163:19:@14249.4]
  wire  storeAddrNotKnownFlags_14_1; // @[LoadQueue.scala 163:19:@14251.4]
  wire  storeAddrNotKnownFlags_14_2; // @[LoadQueue.scala 163:19:@14253.4]
  wire  storeAddrNotKnownFlags_14_3; // @[LoadQueue.scala 163:19:@14255.4]
  wire  storeAddrNotKnownFlags_14_4; // @[LoadQueue.scala 163:19:@14257.4]
  wire  storeAddrNotKnownFlags_14_5; // @[LoadQueue.scala 163:19:@14259.4]
  wire  storeAddrNotKnownFlags_14_6; // @[LoadQueue.scala 163:19:@14261.4]
  wire  storeAddrNotKnownFlags_14_7; // @[LoadQueue.scala 163:19:@14263.4]
  wire  storeAddrNotKnownFlags_14_8; // @[LoadQueue.scala 163:19:@14265.4]
  wire  storeAddrNotKnownFlags_14_9; // @[LoadQueue.scala 163:19:@14267.4]
  wire  storeAddrNotKnownFlags_14_10; // @[LoadQueue.scala 163:19:@14269.4]
  wire  storeAddrNotKnownFlags_14_11; // @[LoadQueue.scala 163:19:@14271.4]
  wire  storeAddrNotKnownFlags_14_12; // @[LoadQueue.scala 163:19:@14273.4]
  wire  storeAddrNotKnownFlags_14_13; // @[LoadQueue.scala 163:19:@14275.4]
  wire  storeAddrNotKnownFlags_14_14; // @[LoadQueue.scala 163:19:@14277.4]
  wire  storeAddrNotKnownFlags_14_15; // @[LoadQueue.scala 163:19:@14279.4]
  wire  storeAddrNotKnownFlags_15_0; // @[LoadQueue.scala 163:19:@14297.4]
  wire  storeAddrNotKnownFlags_15_1; // @[LoadQueue.scala 163:19:@14299.4]
  wire  storeAddrNotKnownFlags_15_2; // @[LoadQueue.scala 163:19:@14301.4]
  wire  storeAddrNotKnownFlags_15_3; // @[LoadQueue.scala 163:19:@14303.4]
  wire  storeAddrNotKnownFlags_15_4; // @[LoadQueue.scala 163:19:@14305.4]
  wire  storeAddrNotKnownFlags_15_5; // @[LoadQueue.scala 163:19:@14307.4]
  wire  storeAddrNotKnownFlags_15_6; // @[LoadQueue.scala 163:19:@14309.4]
  wire  storeAddrNotKnownFlags_15_7; // @[LoadQueue.scala 163:19:@14311.4]
  wire  storeAddrNotKnownFlags_15_8; // @[LoadQueue.scala 163:19:@14313.4]
  wire  storeAddrNotKnownFlags_15_9; // @[LoadQueue.scala 163:19:@14315.4]
  wire  storeAddrNotKnownFlags_15_10; // @[LoadQueue.scala 163:19:@14317.4]
  wire  storeAddrNotKnownFlags_15_11; // @[LoadQueue.scala 163:19:@14319.4]
  wire  storeAddrNotKnownFlags_15_12; // @[LoadQueue.scala 163:19:@14321.4]
  wire  storeAddrNotKnownFlags_15_13; // @[LoadQueue.scala 163:19:@14323.4]
  wire  storeAddrNotKnownFlags_15_14; // @[LoadQueue.scala 163:19:@14325.4]
  wire  storeAddrNotKnownFlags_15_15; // @[LoadQueue.scala 163:19:@14327.4]
  wire [7:0] _T_18010; // @[Mux.scala 19:72:@14658.4]
  wire [7:0] _T_18017; // @[Mux.scala 19:72:@14665.4]
  wire [15:0] _T_18018; // @[Mux.scala 19:72:@14666.4]
  wire [15:0] _T_18020; // @[Mux.scala 19:72:@14667.4]
  wire [7:0] _T_18027; // @[Mux.scala 19:72:@14674.4]
  wire [7:0] _T_18034; // @[Mux.scala 19:72:@14681.4]
  wire [15:0] _T_18035; // @[Mux.scala 19:72:@14682.4]
  wire [15:0] _T_18037; // @[Mux.scala 19:72:@14683.4]
  wire [7:0] _T_18044; // @[Mux.scala 19:72:@14690.4]
  wire [7:0] _T_18051; // @[Mux.scala 19:72:@14697.4]
  wire [15:0] _T_18052; // @[Mux.scala 19:72:@14698.4]
  wire [15:0] _T_18054; // @[Mux.scala 19:72:@14699.4]
  wire [7:0] _T_18061; // @[Mux.scala 19:72:@14706.4]
  wire [7:0] _T_18068; // @[Mux.scala 19:72:@14713.4]
  wire [15:0] _T_18069; // @[Mux.scala 19:72:@14714.4]
  wire [15:0] _T_18071; // @[Mux.scala 19:72:@14715.4]
  wire [7:0] _T_18078; // @[Mux.scala 19:72:@14722.4]
  wire [7:0] _T_18085; // @[Mux.scala 19:72:@14729.4]
  wire [15:0] _T_18086; // @[Mux.scala 19:72:@14730.4]
  wire [15:0] _T_18088; // @[Mux.scala 19:72:@14731.4]
  wire [7:0] _T_18095; // @[Mux.scala 19:72:@14738.4]
  wire [7:0] _T_18102; // @[Mux.scala 19:72:@14745.4]
  wire [15:0] _T_18103; // @[Mux.scala 19:72:@14746.4]
  wire [15:0] _T_18105; // @[Mux.scala 19:72:@14747.4]
  wire [7:0] _T_18112; // @[Mux.scala 19:72:@14754.4]
  wire [7:0] _T_18119; // @[Mux.scala 19:72:@14761.4]
  wire [15:0] _T_18120; // @[Mux.scala 19:72:@14762.4]
  wire [15:0] _T_18122; // @[Mux.scala 19:72:@14763.4]
  wire [7:0] _T_18129; // @[Mux.scala 19:72:@14770.4]
  wire [7:0] _T_18136; // @[Mux.scala 19:72:@14777.4]
  wire [15:0] _T_18137; // @[Mux.scala 19:72:@14778.4]
  wire [15:0] _T_18139; // @[Mux.scala 19:72:@14779.4]
  wire [15:0] _T_18154; // @[Mux.scala 19:72:@14794.4]
  wire [15:0] _T_18156; // @[Mux.scala 19:72:@14795.4]
  wire [15:0] _T_18171; // @[Mux.scala 19:72:@14810.4]
  wire [15:0] _T_18173; // @[Mux.scala 19:72:@14811.4]
  wire [15:0] _T_18188; // @[Mux.scala 19:72:@14826.4]
  wire [15:0] _T_18190; // @[Mux.scala 19:72:@14827.4]
  wire [15:0] _T_18205; // @[Mux.scala 19:72:@14842.4]
  wire [15:0] _T_18207; // @[Mux.scala 19:72:@14843.4]
  wire [15:0] _T_18222; // @[Mux.scala 19:72:@14858.4]
  wire [15:0] _T_18224; // @[Mux.scala 19:72:@14859.4]
  wire [15:0] _T_18239; // @[Mux.scala 19:72:@14874.4]
  wire [15:0] _T_18241; // @[Mux.scala 19:72:@14875.4]
  wire [15:0] _T_18256; // @[Mux.scala 19:72:@14890.4]
  wire [15:0] _T_18258; // @[Mux.scala 19:72:@14891.4]
  wire [15:0] _T_18273; // @[Mux.scala 19:72:@14906.4]
  wire [15:0] _T_18275; // @[Mux.scala 19:72:@14907.4]
  wire [15:0] _T_18276; // @[Mux.scala 19:72:@14908.4]
  wire [15:0] _T_18277; // @[Mux.scala 19:72:@14909.4]
  wire [15:0] _T_18278; // @[Mux.scala 19:72:@14910.4]
  wire [15:0] _T_18279; // @[Mux.scala 19:72:@14911.4]
  wire [15:0] _T_18280; // @[Mux.scala 19:72:@14912.4]
  wire [15:0] _T_18281; // @[Mux.scala 19:72:@14913.4]
  wire [15:0] _T_18282; // @[Mux.scala 19:72:@14914.4]
  wire [15:0] _T_18283; // @[Mux.scala 19:72:@14915.4]
  wire [15:0] _T_18284; // @[Mux.scala 19:72:@14916.4]
  wire [15:0] _T_18285; // @[Mux.scala 19:72:@14917.4]
  wire [15:0] _T_18286; // @[Mux.scala 19:72:@14918.4]
  wire [15:0] _T_18287; // @[Mux.scala 19:72:@14919.4]
  wire [15:0] _T_18288; // @[Mux.scala 19:72:@14920.4]
  wire [15:0] _T_18289; // @[Mux.scala 19:72:@14921.4]
  wire [15:0] _T_18290; // @[Mux.scala 19:72:@14922.4]
  wire [7:0] _T_18868; // @[Mux.scala 19:72:@15272.4]
  wire [7:0] _T_18875; // @[Mux.scala 19:72:@15279.4]
  wire [15:0] _T_18876; // @[Mux.scala 19:72:@15280.4]
  wire [15:0] _T_18878; // @[Mux.scala 19:72:@15281.4]
  wire [7:0] _T_18885; // @[Mux.scala 19:72:@15288.4]
  wire [7:0] _T_18892; // @[Mux.scala 19:72:@15295.4]
  wire [15:0] _T_18893; // @[Mux.scala 19:72:@15296.4]
  wire [15:0] _T_18895; // @[Mux.scala 19:72:@15297.4]
  wire [7:0] _T_18902; // @[Mux.scala 19:72:@15304.4]
  wire [7:0] _T_18909; // @[Mux.scala 19:72:@15311.4]
  wire [15:0] _T_18910; // @[Mux.scala 19:72:@15312.4]
  wire [15:0] _T_18912; // @[Mux.scala 19:72:@15313.4]
  wire [7:0] _T_18919; // @[Mux.scala 19:72:@15320.4]
  wire [7:0] _T_18926; // @[Mux.scala 19:72:@15327.4]
  wire [15:0] _T_18927; // @[Mux.scala 19:72:@15328.4]
  wire [15:0] _T_18929; // @[Mux.scala 19:72:@15329.4]
  wire [7:0] _T_18936; // @[Mux.scala 19:72:@15336.4]
  wire [7:0] _T_18943; // @[Mux.scala 19:72:@15343.4]
  wire [15:0] _T_18944; // @[Mux.scala 19:72:@15344.4]
  wire [15:0] _T_18946; // @[Mux.scala 19:72:@15345.4]
  wire [7:0] _T_18953; // @[Mux.scala 19:72:@15352.4]
  wire [7:0] _T_18960; // @[Mux.scala 19:72:@15359.4]
  wire [15:0] _T_18961; // @[Mux.scala 19:72:@15360.4]
  wire [15:0] _T_18963; // @[Mux.scala 19:72:@15361.4]
  wire [7:0] _T_18970; // @[Mux.scala 19:72:@15368.4]
  wire [7:0] _T_18977; // @[Mux.scala 19:72:@15375.4]
  wire [15:0] _T_18978; // @[Mux.scala 19:72:@15376.4]
  wire [15:0] _T_18980; // @[Mux.scala 19:72:@15377.4]
  wire [7:0] _T_18987; // @[Mux.scala 19:72:@15384.4]
  wire [7:0] _T_18994; // @[Mux.scala 19:72:@15391.4]
  wire [15:0] _T_18995; // @[Mux.scala 19:72:@15392.4]
  wire [15:0] _T_18997; // @[Mux.scala 19:72:@15393.4]
  wire [15:0] _T_19012; // @[Mux.scala 19:72:@15408.4]
  wire [15:0] _T_19014; // @[Mux.scala 19:72:@15409.4]
  wire [15:0] _T_19029; // @[Mux.scala 19:72:@15424.4]
  wire [15:0] _T_19031; // @[Mux.scala 19:72:@15425.4]
  wire [15:0] _T_19046; // @[Mux.scala 19:72:@15440.4]
  wire [15:0] _T_19048; // @[Mux.scala 19:72:@15441.4]
  wire [15:0] _T_19063; // @[Mux.scala 19:72:@15456.4]
  wire [15:0] _T_19065; // @[Mux.scala 19:72:@15457.4]
  wire [15:0] _T_19080; // @[Mux.scala 19:72:@15472.4]
  wire [15:0] _T_19082; // @[Mux.scala 19:72:@15473.4]
  wire [15:0] _T_19097; // @[Mux.scala 19:72:@15488.4]
  wire [15:0] _T_19099; // @[Mux.scala 19:72:@15489.4]
  wire [15:0] _T_19114; // @[Mux.scala 19:72:@15504.4]
  wire [15:0] _T_19116; // @[Mux.scala 19:72:@15505.4]
  wire [15:0] _T_19131; // @[Mux.scala 19:72:@15520.4]
  wire [15:0] _T_19133; // @[Mux.scala 19:72:@15521.4]
  wire [15:0] _T_19134; // @[Mux.scala 19:72:@15522.4]
  wire [15:0] _T_19135; // @[Mux.scala 19:72:@15523.4]
  wire [15:0] _T_19136; // @[Mux.scala 19:72:@15524.4]
  wire [15:0] _T_19137; // @[Mux.scala 19:72:@15525.4]
  wire [15:0] _T_19138; // @[Mux.scala 19:72:@15526.4]
  wire [15:0] _T_19139; // @[Mux.scala 19:72:@15527.4]
  wire [15:0] _T_19140; // @[Mux.scala 19:72:@15528.4]
  wire [15:0] _T_19141; // @[Mux.scala 19:72:@15529.4]
  wire [15:0] _T_19142; // @[Mux.scala 19:72:@15530.4]
  wire [15:0] _T_19143; // @[Mux.scala 19:72:@15531.4]
  wire [15:0] _T_19144; // @[Mux.scala 19:72:@15532.4]
  wire [15:0] _T_19145; // @[Mux.scala 19:72:@15533.4]
  wire [15:0] _T_19146; // @[Mux.scala 19:72:@15534.4]
  wire [15:0] _T_19147; // @[Mux.scala 19:72:@15535.4]
  wire [15:0] _T_19148; // @[Mux.scala 19:72:@15536.4]
  wire [7:0] _T_19726; // @[Mux.scala 19:72:@15886.4]
  wire [7:0] _T_19733; // @[Mux.scala 19:72:@15893.4]
  wire [15:0] _T_19734; // @[Mux.scala 19:72:@15894.4]
  wire [15:0] _T_19736; // @[Mux.scala 19:72:@15895.4]
  wire [7:0] _T_19743; // @[Mux.scala 19:72:@15902.4]
  wire [7:0] _T_19750; // @[Mux.scala 19:72:@15909.4]
  wire [15:0] _T_19751; // @[Mux.scala 19:72:@15910.4]
  wire [15:0] _T_19753; // @[Mux.scala 19:72:@15911.4]
  wire [7:0] _T_19760; // @[Mux.scala 19:72:@15918.4]
  wire [7:0] _T_19767; // @[Mux.scala 19:72:@15925.4]
  wire [15:0] _T_19768; // @[Mux.scala 19:72:@15926.4]
  wire [15:0] _T_19770; // @[Mux.scala 19:72:@15927.4]
  wire [7:0] _T_19777; // @[Mux.scala 19:72:@15934.4]
  wire [7:0] _T_19784; // @[Mux.scala 19:72:@15941.4]
  wire [15:0] _T_19785; // @[Mux.scala 19:72:@15942.4]
  wire [15:0] _T_19787; // @[Mux.scala 19:72:@15943.4]
  wire [7:0] _T_19794; // @[Mux.scala 19:72:@15950.4]
  wire [7:0] _T_19801; // @[Mux.scala 19:72:@15957.4]
  wire [15:0] _T_19802; // @[Mux.scala 19:72:@15958.4]
  wire [15:0] _T_19804; // @[Mux.scala 19:72:@15959.4]
  wire [7:0] _T_19811; // @[Mux.scala 19:72:@15966.4]
  wire [7:0] _T_19818; // @[Mux.scala 19:72:@15973.4]
  wire [15:0] _T_19819; // @[Mux.scala 19:72:@15974.4]
  wire [15:0] _T_19821; // @[Mux.scala 19:72:@15975.4]
  wire [7:0] _T_19828; // @[Mux.scala 19:72:@15982.4]
  wire [7:0] _T_19835; // @[Mux.scala 19:72:@15989.4]
  wire [15:0] _T_19836; // @[Mux.scala 19:72:@15990.4]
  wire [15:0] _T_19838; // @[Mux.scala 19:72:@15991.4]
  wire [7:0] _T_19845; // @[Mux.scala 19:72:@15998.4]
  wire [7:0] _T_19852; // @[Mux.scala 19:72:@16005.4]
  wire [15:0] _T_19853; // @[Mux.scala 19:72:@16006.4]
  wire [15:0] _T_19855; // @[Mux.scala 19:72:@16007.4]
  wire [15:0] _T_19870; // @[Mux.scala 19:72:@16022.4]
  wire [15:0] _T_19872; // @[Mux.scala 19:72:@16023.4]
  wire [15:0] _T_19887; // @[Mux.scala 19:72:@16038.4]
  wire [15:0] _T_19889; // @[Mux.scala 19:72:@16039.4]
  wire [15:0] _T_19904; // @[Mux.scala 19:72:@16054.4]
  wire [15:0] _T_19906; // @[Mux.scala 19:72:@16055.4]
  wire [15:0] _T_19921; // @[Mux.scala 19:72:@16070.4]
  wire [15:0] _T_19923; // @[Mux.scala 19:72:@16071.4]
  wire [15:0] _T_19938; // @[Mux.scala 19:72:@16086.4]
  wire [15:0] _T_19940; // @[Mux.scala 19:72:@16087.4]
  wire [15:0] _T_19955; // @[Mux.scala 19:72:@16102.4]
  wire [15:0] _T_19957; // @[Mux.scala 19:72:@16103.4]
  wire [15:0] _T_19972; // @[Mux.scala 19:72:@16118.4]
  wire [15:0] _T_19974; // @[Mux.scala 19:72:@16119.4]
  wire [15:0] _T_19989; // @[Mux.scala 19:72:@16134.4]
  wire [15:0] _T_19991; // @[Mux.scala 19:72:@16135.4]
  wire [15:0] _T_19992; // @[Mux.scala 19:72:@16136.4]
  wire [15:0] _T_19993; // @[Mux.scala 19:72:@16137.4]
  wire [15:0] _T_19994; // @[Mux.scala 19:72:@16138.4]
  wire [15:0] _T_19995; // @[Mux.scala 19:72:@16139.4]
  wire [15:0] _T_19996; // @[Mux.scala 19:72:@16140.4]
  wire [15:0] _T_19997; // @[Mux.scala 19:72:@16141.4]
  wire [15:0] _T_19998; // @[Mux.scala 19:72:@16142.4]
  wire [15:0] _T_19999; // @[Mux.scala 19:72:@16143.4]
  wire [15:0] _T_20000; // @[Mux.scala 19:72:@16144.4]
  wire [15:0] _T_20001; // @[Mux.scala 19:72:@16145.4]
  wire [15:0] _T_20002; // @[Mux.scala 19:72:@16146.4]
  wire [15:0] _T_20003; // @[Mux.scala 19:72:@16147.4]
  wire [15:0] _T_20004; // @[Mux.scala 19:72:@16148.4]
  wire [15:0] _T_20005; // @[Mux.scala 19:72:@16149.4]
  wire [15:0] _T_20006; // @[Mux.scala 19:72:@16150.4]
  wire [7:0] _T_20584; // @[Mux.scala 19:72:@16500.4]
  wire [7:0] _T_20591; // @[Mux.scala 19:72:@16507.4]
  wire [15:0] _T_20592; // @[Mux.scala 19:72:@16508.4]
  wire [15:0] _T_20594; // @[Mux.scala 19:72:@16509.4]
  wire [7:0] _T_20601; // @[Mux.scala 19:72:@16516.4]
  wire [7:0] _T_20608; // @[Mux.scala 19:72:@16523.4]
  wire [15:0] _T_20609; // @[Mux.scala 19:72:@16524.4]
  wire [15:0] _T_20611; // @[Mux.scala 19:72:@16525.4]
  wire [7:0] _T_20618; // @[Mux.scala 19:72:@16532.4]
  wire [7:0] _T_20625; // @[Mux.scala 19:72:@16539.4]
  wire [15:0] _T_20626; // @[Mux.scala 19:72:@16540.4]
  wire [15:0] _T_20628; // @[Mux.scala 19:72:@16541.4]
  wire [7:0] _T_20635; // @[Mux.scala 19:72:@16548.4]
  wire [7:0] _T_20642; // @[Mux.scala 19:72:@16555.4]
  wire [15:0] _T_20643; // @[Mux.scala 19:72:@16556.4]
  wire [15:0] _T_20645; // @[Mux.scala 19:72:@16557.4]
  wire [7:0] _T_20652; // @[Mux.scala 19:72:@16564.4]
  wire [7:0] _T_20659; // @[Mux.scala 19:72:@16571.4]
  wire [15:0] _T_20660; // @[Mux.scala 19:72:@16572.4]
  wire [15:0] _T_20662; // @[Mux.scala 19:72:@16573.4]
  wire [7:0] _T_20669; // @[Mux.scala 19:72:@16580.4]
  wire [7:0] _T_20676; // @[Mux.scala 19:72:@16587.4]
  wire [15:0] _T_20677; // @[Mux.scala 19:72:@16588.4]
  wire [15:0] _T_20679; // @[Mux.scala 19:72:@16589.4]
  wire [7:0] _T_20686; // @[Mux.scala 19:72:@16596.4]
  wire [7:0] _T_20693; // @[Mux.scala 19:72:@16603.4]
  wire [15:0] _T_20694; // @[Mux.scala 19:72:@16604.4]
  wire [15:0] _T_20696; // @[Mux.scala 19:72:@16605.4]
  wire [7:0] _T_20703; // @[Mux.scala 19:72:@16612.4]
  wire [7:0] _T_20710; // @[Mux.scala 19:72:@16619.4]
  wire [15:0] _T_20711; // @[Mux.scala 19:72:@16620.4]
  wire [15:0] _T_20713; // @[Mux.scala 19:72:@16621.4]
  wire [15:0] _T_20728; // @[Mux.scala 19:72:@16636.4]
  wire [15:0] _T_20730; // @[Mux.scala 19:72:@16637.4]
  wire [15:0] _T_20745; // @[Mux.scala 19:72:@16652.4]
  wire [15:0] _T_20747; // @[Mux.scala 19:72:@16653.4]
  wire [15:0] _T_20762; // @[Mux.scala 19:72:@16668.4]
  wire [15:0] _T_20764; // @[Mux.scala 19:72:@16669.4]
  wire [15:0] _T_20779; // @[Mux.scala 19:72:@16684.4]
  wire [15:0] _T_20781; // @[Mux.scala 19:72:@16685.4]
  wire [15:0] _T_20796; // @[Mux.scala 19:72:@16700.4]
  wire [15:0] _T_20798; // @[Mux.scala 19:72:@16701.4]
  wire [15:0] _T_20813; // @[Mux.scala 19:72:@16716.4]
  wire [15:0] _T_20815; // @[Mux.scala 19:72:@16717.4]
  wire [15:0] _T_20830; // @[Mux.scala 19:72:@16732.4]
  wire [15:0] _T_20832; // @[Mux.scala 19:72:@16733.4]
  wire [15:0] _T_20847; // @[Mux.scala 19:72:@16748.4]
  wire [15:0] _T_20849; // @[Mux.scala 19:72:@16749.4]
  wire [15:0] _T_20850; // @[Mux.scala 19:72:@16750.4]
  wire [15:0] _T_20851; // @[Mux.scala 19:72:@16751.4]
  wire [15:0] _T_20852; // @[Mux.scala 19:72:@16752.4]
  wire [15:0] _T_20853; // @[Mux.scala 19:72:@16753.4]
  wire [15:0] _T_20854; // @[Mux.scala 19:72:@16754.4]
  wire [15:0] _T_20855; // @[Mux.scala 19:72:@16755.4]
  wire [15:0] _T_20856; // @[Mux.scala 19:72:@16756.4]
  wire [15:0] _T_20857; // @[Mux.scala 19:72:@16757.4]
  wire [15:0] _T_20858; // @[Mux.scala 19:72:@16758.4]
  wire [15:0] _T_20859; // @[Mux.scala 19:72:@16759.4]
  wire [15:0] _T_20860; // @[Mux.scala 19:72:@16760.4]
  wire [15:0] _T_20861; // @[Mux.scala 19:72:@16761.4]
  wire [15:0] _T_20862; // @[Mux.scala 19:72:@16762.4]
  wire [15:0] _T_20863; // @[Mux.scala 19:72:@16763.4]
  wire [15:0] _T_20864; // @[Mux.scala 19:72:@16764.4]
  wire [7:0] _T_21442; // @[Mux.scala 19:72:@17114.4]
  wire [7:0] _T_21449; // @[Mux.scala 19:72:@17121.4]
  wire [15:0] _T_21450; // @[Mux.scala 19:72:@17122.4]
  wire [15:0] _T_21452; // @[Mux.scala 19:72:@17123.4]
  wire [7:0] _T_21459; // @[Mux.scala 19:72:@17130.4]
  wire [7:0] _T_21466; // @[Mux.scala 19:72:@17137.4]
  wire [15:0] _T_21467; // @[Mux.scala 19:72:@17138.4]
  wire [15:0] _T_21469; // @[Mux.scala 19:72:@17139.4]
  wire [7:0] _T_21476; // @[Mux.scala 19:72:@17146.4]
  wire [7:0] _T_21483; // @[Mux.scala 19:72:@17153.4]
  wire [15:0] _T_21484; // @[Mux.scala 19:72:@17154.4]
  wire [15:0] _T_21486; // @[Mux.scala 19:72:@17155.4]
  wire [7:0] _T_21493; // @[Mux.scala 19:72:@17162.4]
  wire [7:0] _T_21500; // @[Mux.scala 19:72:@17169.4]
  wire [15:0] _T_21501; // @[Mux.scala 19:72:@17170.4]
  wire [15:0] _T_21503; // @[Mux.scala 19:72:@17171.4]
  wire [7:0] _T_21510; // @[Mux.scala 19:72:@17178.4]
  wire [7:0] _T_21517; // @[Mux.scala 19:72:@17185.4]
  wire [15:0] _T_21518; // @[Mux.scala 19:72:@17186.4]
  wire [15:0] _T_21520; // @[Mux.scala 19:72:@17187.4]
  wire [7:0] _T_21527; // @[Mux.scala 19:72:@17194.4]
  wire [7:0] _T_21534; // @[Mux.scala 19:72:@17201.4]
  wire [15:0] _T_21535; // @[Mux.scala 19:72:@17202.4]
  wire [15:0] _T_21537; // @[Mux.scala 19:72:@17203.4]
  wire [7:0] _T_21544; // @[Mux.scala 19:72:@17210.4]
  wire [7:0] _T_21551; // @[Mux.scala 19:72:@17217.4]
  wire [15:0] _T_21552; // @[Mux.scala 19:72:@17218.4]
  wire [15:0] _T_21554; // @[Mux.scala 19:72:@17219.4]
  wire [7:0] _T_21561; // @[Mux.scala 19:72:@17226.4]
  wire [7:0] _T_21568; // @[Mux.scala 19:72:@17233.4]
  wire [15:0] _T_21569; // @[Mux.scala 19:72:@17234.4]
  wire [15:0] _T_21571; // @[Mux.scala 19:72:@17235.4]
  wire [15:0] _T_21586; // @[Mux.scala 19:72:@17250.4]
  wire [15:0] _T_21588; // @[Mux.scala 19:72:@17251.4]
  wire [15:0] _T_21603; // @[Mux.scala 19:72:@17266.4]
  wire [15:0] _T_21605; // @[Mux.scala 19:72:@17267.4]
  wire [15:0] _T_21620; // @[Mux.scala 19:72:@17282.4]
  wire [15:0] _T_21622; // @[Mux.scala 19:72:@17283.4]
  wire [15:0] _T_21637; // @[Mux.scala 19:72:@17298.4]
  wire [15:0] _T_21639; // @[Mux.scala 19:72:@17299.4]
  wire [15:0] _T_21654; // @[Mux.scala 19:72:@17314.4]
  wire [15:0] _T_21656; // @[Mux.scala 19:72:@17315.4]
  wire [15:0] _T_21671; // @[Mux.scala 19:72:@17330.4]
  wire [15:0] _T_21673; // @[Mux.scala 19:72:@17331.4]
  wire [15:0] _T_21688; // @[Mux.scala 19:72:@17346.4]
  wire [15:0] _T_21690; // @[Mux.scala 19:72:@17347.4]
  wire [15:0] _T_21705; // @[Mux.scala 19:72:@17362.4]
  wire [15:0] _T_21707; // @[Mux.scala 19:72:@17363.4]
  wire [15:0] _T_21708; // @[Mux.scala 19:72:@17364.4]
  wire [15:0] _T_21709; // @[Mux.scala 19:72:@17365.4]
  wire [15:0] _T_21710; // @[Mux.scala 19:72:@17366.4]
  wire [15:0] _T_21711; // @[Mux.scala 19:72:@17367.4]
  wire [15:0] _T_21712; // @[Mux.scala 19:72:@17368.4]
  wire [15:0] _T_21713; // @[Mux.scala 19:72:@17369.4]
  wire [15:0] _T_21714; // @[Mux.scala 19:72:@17370.4]
  wire [15:0] _T_21715; // @[Mux.scala 19:72:@17371.4]
  wire [15:0] _T_21716; // @[Mux.scala 19:72:@17372.4]
  wire [15:0] _T_21717; // @[Mux.scala 19:72:@17373.4]
  wire [15:0] _T_21718; // @[Mux.scala 19:72:@17374.4]
  wire [15:0] _T_21719; // @[Mux.scala 19:72:@17375.4]
  wire [15:0] _T_21720; // @[Mux.scala 19:72:@17376.4]
  wire [15:0] _T_21721; // @[Mux.scala 19:72:@17377.4]
  wire [15:0] _T_21722; // @[Mux.scala 19:72:@17378.4]
  wire [7:0] _T_22300; // @[Mux.scala 19:72:@17728.4]
  wire [7:0] _T_22307; // @[Mux.scala 19:72:@17735.4]
  wire [15:0] _T_22308; // @[Mux.scala 19:72:@17736.4]
  wire [15:0] _T_22310; // @[Mux.scala 19:72:@17737.4]
  wire [7:0] _T_22317; // @[Mux.scala 19:72:@17744.4]
  wire [7:0] _T_22324; // @[Mux.scala 19:72:@17751.4]
  wire [15:0] _T_22325; // @[Mux.scala 19:72:@17752.4]
  wire [15:0] _T_22327; // @[Mux.scala 19:72:@17753.4]
  wire [7:0] _T_22334; // @[Mux.scala 19:72:@17760.4]
  wire [7:0] _T_22341; // @[Mux.scala 19:72:@17767.4]
  wire [15:0] _T_22342; // @[Mux.scala 19:72:@17768.4]
  wire [15:0] _T_22344; // @[Mux.scala 19:72:@17769.4]
  wire [7:0] _T_22351; // @[Mux.scala 19:72:@17776.4]
  wire [7:0] _T_22358; // @[Mux.scala 19:72:@17783.4]
  wire [15:0] _T_22359; // @[Mux.scala 19:72:@17784.4]
  wire [15:0] _T_22361; // @[Mux.scala 19:72:@17785.4]
  wire [7:0] _T_22368; // @[Mux.scala 19:72:@17792.4]
  wire [7:0] _T_22375; // @[Mux.scala 19:72:@17799.4]
  wire [15:0] _T_22376; // @[Mux.scala 19:72:@17800.4]
  wire [15:0] _T_22378; // @[Mux.scala 19:72:@17801.4]
  wire [7:0] _T_22385; // @[Mux.scala 19:72:@17808.4]
  wire [7:0] _T_22392; // @[Mux.scala 19:72:@17815.4]
  wire [15:0] _T_22393; // @[Mux.scala 19:72:@17816.4]
  wire [15:0] _T_22395; // @[Mux.scala 19:72:@17817.4]
  wire [7:0] _T_22402; // @[Mux.scala 19:72:@17824.4]
  wire [7:0] _T_22409; // @[Mux.scala 19:72:@17831.4]
  wire [15:0] _T_22410; // @[Mux.scala 19:72:@17832.4]
  wire [15:0] _T_22412; // @[Mux.scala 19:72:@17833.4]
  wire [7:0] _T_22419; // @[Mux.scala 19:72:@17840.4]
  wire [7:0] _T_22426; // @[Mux.scala 19:72:@17847.4]
  wire [15:0] _T_22427; // @[Mux.scala 19:72:@17848.4]
  wire [15:0] _T_22429; // @[Mux.scala 19:72:@17849.4]
  wire [15:0] _T_22444; // @[Mux.scala 19:72:@17864.4]
  wire [15:0] _T_22446; // @[Mux.scala 19:72:@17865.4]
  wire [15:0] _T_22461; // @[Mux.scala 19:72:@17880.4]
  wire [15:0] _T_22463; // @[Mux.scala 19:72:@17881.4]
  wire [15:0] _T_22478; // @[Mux.scala 19:72:@17896.4]
  wire [15:0] _T_22480; // @[Mux.scala 19:72:@17897.4]
  wire [15:0] _T_22495; // @[Mux.scala 19:72:@17912.4]
  wire [15:0] _T_22497; // @[Mux.scala 19:72:@17913.4]
  wire [15:0] _T_22512; // @[Mux.scala 19:72:@17928.4]
  wire [15:0] _T_22514; // @[Mux.scala 19:72:@17929.4]
  wire [15:0] _T_22529; // @[Mux.scala 19:72:@17944.4]
  wire [15:0] _T_22531; // @[Mux.scala 19:72:@17945.4]
  wire [15:0] _T_22546; // @[Mux.scala 19:72:@17960.4]
  wire [15:0] _T_22548; // @[Mux.scala 19:72:@17961.4]
  wire [15:0] _T_22563; // @[Mux.scala 19:72:@17976.4]
  wire [15:0] _T_22565; // @[Mux.scala 19:72:@17977.4]
  wire [15:0] _T_22566; // @[Mux.scala 19:72:@17978.4]
  wire [15:0] _T_22567; // @[Mux.scala 19:72:@17979.4]
  wire [15:0] _T_22568; // @[Mux.scala 19:72:@17980.4]
  wire [15:0] _T_22569; // @[Mux.scala 19:72:@17981.4]
  wire [15:0] _T_22570; // @[Mux.scala 19:72:@17982.4]
  wire [15:0] _T_22571; // @[Mux.scala 19:72:@17983.4]
  wire [15:0] _T_22572; // @[Mux.scala 19:72:@17984.4]
  wire [15:0] _T_22573; // @[Mux.scala 19:72:@17985.4]
  wire [15:0] _T_22574; // @[Mux.scala 19:72:@17986.4]
  wire [15:0] _T_22575; // @[Mux.scala 19:72:@17987.4]
  wire [15:0] _T_22576; // @[Mux.scala 19:72:@17988.4]
  wire [15:0] _T_22577; // @[Mux.scala 19:72:@17989.4]
  wire [15:0] _T_22578; // @[Mux.scala 19:72:@17990.4]
  wire [15:0] _T_22579; // @[Mux.scala 19:72:@17991.4]
  wire [15:0] _T_22580; // @[Mux.scala 19:72:@17992.4]
  wire [7:0] _T_23158; // @[Mux.scala 19:72:@18342.4]
  wire [7:0] _T_23165; // @[Mux.scala 19:72:@18349.4]
  wire [15:0] _T_23166; // @[Mux.scala 19:72:@18350.4]
  wire [15:0] _T_23168; // @[Mux.scala 19:72:@18351.4]
  wire [7:0] _T_23175; // @[Mux.scala 19:72:@18358.4]
  wire [7:0] _T_23182; // @[Mux.scala 19:72:@18365.4]
  wire [15:0] _T_23183; // @[Mux.scala 19:72:@18366.4]
  wire [15:0] _T_23185; // @[Mux.scala 19:72:@18367.4]
  wire [7:0] _T_23192; // @[Mux.scala 19:72:@18374.4]
  wire [7:0] _T_23199; // @[Mux.scala 19:72:@18381.4]
  wire [15:0] _T_23200; // @[Mux.scala 19:72:@18382.4]
  wire [15:0] _T_23202; // @[Mux.scala 19:72:@18383.4]
  wire [7:0] _T_23209; // @[Mux.scala 19:72:@18390.4]
  wire [7:0] _T_23216; // @[Mux.scala 19:72:@18397.4]
  wire [15:0] _T_23217; // @[Mux.scala 19:72:@18398.4]
  wire [15:0] _T_23219; // @[Mux.scala 19:72:@18399.4]
  wire [7:0] _T_23226; // @[Mux.scala 19:72:@18406.4]
  wire [7:0] _T_23233; // @[Mux.scala 19:72:@18413.4]
  wire [15:0] _T_23234; // @[Mux.scala 19:72:@18414.4]
  wire [15:0] _T_23236; // @[Mux.scala 19:72:@18415.4]
  wire [7:0] _T_23243; // @[Mux.scala 19:72:@18422.4]
  wire [7:0] _T_23250; // @[Mux.scala 19:72:@18429.4]
  wire [15:0] _T_23251; // @[Mux.scala 19:72:@18430.4]
  wire [15:0] _T_23253; // @[Mux.scala 19:72:@18431.4]
  wire [7:0] _T_23260; // @[Mux.scala 19:72:@18438.4]
  wire [7:0] _T_23267; // @[Mux.scala 19:72:@18445.4]
  wire [15:0] _T_23268; // @[Mux.scala 19:72:@18446.4]
  wire [15:0] _T_23270; // @[Mux.scala 19:72:@18447.4]
  wire [7:0] _T_23277; // @[Mux.scala 19:72:@18454.4]
  wire [7:0] _T_23284; // @[Mux.scala 19:72:@18461.4]
  wire [15:0] _T_23285; // @[Mux.scala 19:72:@18462.4]
  wire [15:0] _T_23287; // @[Mux.scala 19:72:@18463.4]
  wire [15:0] _T_23302; // @[Mux.scala 19:72:@18478.4]
  wire [15:0] _T_23304; // @[Mux.scala 19:72:@18479.4]
  wire [15:0] _T_23319; // @[Mux.scala 19:72:@18494.4]
  wire [15:0] _T_23321; // @[Mux.scala 19:72:@18495.4]
  wire [15:0] _T_23336; // @[Mux.scala 19:72:@18510.4]
  wire [15:0] _T_23338; // @[Mux.scala 19:72:@18511.4]
  wire [15:0] _T_23353; // @[Mux.scala 19:72:@18526.4]
  wire [15:0] _T_23355; // @[Mux.scala 19:72:@18527.4]
  wire [15:0] _T_23370; // @[Mux.scala 19:72:@18542.4]
  wire [15:0] _T_23372; // @[Mux.scala 19:72:@18543.4]
  wire [15:0] _T_23387; // @[Mux.scala 19:72:@18558.4]
  wire [15:0] _T_23389; // @[Mux.scala 19:72:@18559.4]
  wire [15:0] _T_23404; // @[Mux.scala 19:72:@18574.4]
  wire [15:0] _T_23406; // @[Mux.scala 19:72:@18575.4]
  wire [15:0] _T_23421; // @[Mux.scala 19:72:@18590.4]
  wire [15:0] _T_23423; // @[Mux.scala 19:72:@18591.4]
  wire [15:0] _T_23424; // @[Mux.scala 19:72:@18592.4]
  wire [15:0] _T_23425; // @[Mux.scala 19:72:@18593.4]
  wire [15:0] _T_23426; // @[Mux.scala 19:72:@18594.4]
  wire [15:0] _T_23427; // @[Mux.scala 19:72:@18595.4]
  wire [15:0] _T_23428; // @[Mux.scala 19:72:@18596.4]
  wire [15:0] _T_23429; // @[Mux.scala 19:72:@18597.4]
  wire [15:0] _T_23430; // @[Mux.scala 19:72:@18598.4]
  wire [15:0] _T_23431; // @[Mux.scala 19:72:@18599.4]
  wire [15:0] _T_23432; // @[Mux.scala 19:72:@18600.4]
  wire [15:0] _T_23433; // @[Mux.scala 19:72:@18601.4]
  wire [15:0] _T_23434; // @[Mux.scala 19:72:@18602.4]
  wire [15:0] _T_23435; // @[Mux.scala 19:72:@18603.4]
  wire [15:0] _T_23436; // @[Mux.scala 19:72:@18604.4]
  wire [15:0] _T_23437; // @[Mux.scala 19:72:@18605.4]
  wire [15:0] _T_23438; // @[Mux.scala 19:72:@18606.4]
  wire [7:0] _T_24016; // @[Mux.scala 19:72:@18956.4]
  wire [7:0] _T_24023; // @[Mux.scala 19:72:@18963.4]
  wire [15:0] _T_24024; // @[Mux.scala 19:72:@18964.4]
  wire [15:0] _T_24026; // @[Mux.scala 19:72:@18965.4]
  wire [7:0] _T_24033; // @[Mux.scala 19:72:@18972.4]
  wire [7:0] _T_24040; // @[Mux.scala 19:72:@18979.4]
  wire [15:0] _T_24041; // @[Mux.scala 19:72:@18980.4]
  wire [15:0] _T_24043; // @[Mux.scala 19:72:@18981.4]
  wire [7:0] _T_24050; // @[Mux.scala 19:72:@18988.4]
  wire [7:0] _T_24057; // @[Mux.scala 19:72:@18995.4]
  wire [15:0] _T_24058; // @[Mux.scala 19:72:@18996.4]
  wire [15:0] _T_24060; // @[Mux.scala 19:72:@18997.4]
  wire [7:0] _T_24067; // @[Mux.scala 19:72:@19004.4]
  wire [7:0] _T_24074; // @[Mux.scala 19:72:@19011.4]
  wire [15:0] _T_24075; // @[Mux.scala 19:72:@19012.4]
  wire [15:0] _T_24077; // @[Mux.scala 19:72:@19013.4]
  wire [7:0] _T_24084; // @[Mux.scala 19:72:@19020.4]
  wire [7:0] _T_24091; // @[Mux.scala 19:72:@19027.4]
  wire [15:0] _T_24092; // @[Mux.scala 19:72:@19028.4]
  wire [15:0] _T_24094; // @[Mux.scala 19:72:@19029.4]
  wire [7:0] _T_24101; // @[Mux.scala 19:72:@19036.4]
  wire [7:0] _T_24108; // @[Mux.scala 19:72:@19043.4]
  wire [15:0] _T_24109; // @[Mux.scala 19:72:@19044.4]
  wire [15:0] _T_24111; // @[Mux.scala 19:72:@19045.4]
  wire [7:0] _T_24118; // @[Mux.scala 19:72:@19052.4]
  wire [7:0] _T_24125; // @[Mux.scala 19:72:@19059.4]
  wire [15:0] _T_24126; // @[Mux.scala 19:72:@19060.4]
  wire [15:0] _T_24128; // @[Mux.scala 19:72:@19061.4]
  wire [7:0] _T_24135; // @[Mux.scala 19:72:@19068.4]
  wire [7:0] _T_24142; // @[Mux.scala 19:72:@19075.4]
  wire [15:0] _T_24143; // @[Mux.scala 19:72:@19076.4]
  wire [15:0] _T_24145; // @[Mux.scala 19:72:@19077.4]
  wire [15:0] _T_24160; // @[Mux.scala 19:72:@19092.4]
  wire [15:0] _T_24162; // @[Mux.scala 19:72:@19093.4]
  wire [15:0] _T_24177; // @[Mux.scala 19:72:@19108.4]
  wire [15:0] _T_24179; // @[Mux.scala 19:72:@19109.4]
  wire [15:0] _T_24194; // @[Mux.scala 19:72:@19124.4]
  wire [15:0] _T_24196; // @[Mux.scala 19:72:@19125.4]
  wire [15:0] _T_24211; // @[Mux.scala 19:72:@19140.4]
  wire [15:0] _T_24213; // @[Mux.scala 19:72:@19141.4]
  wire [15:0] _T_24228; // @[Mux.scala 19:72:@19156.4]
  wire [15:0] _T_24230; // @[Mux.scala 19:72:@19157.4]
  wire [15:0] _T_24245; // @[Mux.scala 19:72:@19172.4]
  wire [15:0] _T_24247; // @[Mux.scala 19:72:@19173.4]
  wire [15:0] _T_24262; // @[Mux.scala 19:72:@19188.4]
  wire [15:0] _T_24264; // @[Mux.scala 19:72:@19189.4]
  wire [15:0] _T_24279; // @[Mux.scala 19:72:@19204.4]
  wire [15:0] _T_24281; // @[Mux.scala 19:72:@19205.4]
  wire [15:0] _T_24282; // @[Mux.scala 19:72:@19206.4]
  wire [15:0] _T_24283; // @[Mux.scala 19:72:@19207.4]
  wire [15:0] _T_24284; // @[Mux.scala 19:72:@19208.4]
  wire [15:0] _T_24285; // @[Mux.scala 19:72:@19209.4]
  wire [15:0] _T_24286; // @[Mux.scala 19:72:@19210.4]
  wire [15:0] _T_24287; // @[Mux.scala 19:72:@19211.4]
  wire [15:0] _T_24288; // @[Mux.scala 19:72:@19212.4]
  wire [15:0] _T_24289; // @[Mux.scala 19:72:@19213.4]
  wire [15:0] _T_24290; // @[Mux.scala 19:72:@19214.4]
  wire [15:0] _T_24291; // @[Mux.scala 19:72:@19215.4]
  wire [15:0] _T_24292; // @[Mux.scala 19:72:@19216.4]
  wire [15:0] _T_24293; // @[Mux.scala 19:72:@19217.4]
  wire [15:0] _T_24294; // @[Mux.scala 19:72:@19218.4]
  wire [15:0] _T_24295; // @[Mux.scala 19:72:@19219.4]
  wire [15:0] _T_24296; // @[Mux.scala 19:72:@19220.4]
  wire [7:0] _T_24874; // @[Mux.scala 19:72:@19570.4]
  wire [7:0] _T_24881; // @[Mux.scala 19:72:@19577.4]
  wire [15:0] _T_24882; // @[Mux.scala 19:72:@19578.4]
  wire [15:0] _T_24884; // @[Mux.scala 19:72:@19579.4]
  wire [7:0] _T_24891; // @[Mux.scala 19:72:@19586.4]
  wire [7:0] _T_24898; // @[Mux.scala 19:72:@19593.4]
  wire [15:0] _T_24899; // @[Mux.scala 19:72:@19594.4]
  wire [15:0] _T_24901; // @[Mux.scala 19:72:@19595.4]
  wire [7:0] _T_24908; // @[Mux.scala 19:72:@19602.4]
  wire [7:0] _T_24915; // @[Mux.scala 19:72:@19609.4]
  wire [15:0] _T_24916; // @[Mux.scala 19:72:@19610.4]
  wire [15:0] _T_24918; // @[Mux.scala 19:72:@19611.4]
  wire [7:0] _T_24925; // @[Mux.scala 19:72:@19618.4]
  wire [7:0] _T_24932; // @[Mux.scala 19:72:@19625.4]
  wire [15:0] _T_24933; // @[Mux.scala 19:72:@19626.4]
  wire [15:0] _T_24935; // @[Mux.scala 19:72:@19627.4]
  wire [7:0] _T_24942; // @[Mux.scala 19:72:@19634.4]
  wire [7:0] _T_24949; // @[Mux.scala 19:72:@19641.4]
  wire [15:0] _T_24950; // @[Mux.scala 19:72:@19642.4]
  wire [15:0] _T_24952; // @[Mux.scala 19:72:@19643.4]
  wire [7:0] _T_24959; // @[Mux.scala 19:72:@19650.4]
  wire [7:0] _T_24966; // @[Mux.scala 19:72:@19657.4]
  wire [15:0] _T_24967; // @[Mux.scala 19:72:@19658.4]
  wire [15:0] _T_24969; // @[Mux.scala 19:72:@19659.4]
  wire [7:0] _T_24976; // @[Mux.scala 19:72:@19666.4]
  wire [7:0] _T_24983; // @[Mux.scala 19:72:@19673.4]
  wire [15:0] _T_24984; // @[Mux.scala 19:72:@19674.4]
  wire [15:0] _T_24986; // @[Mux.scala 19:72:@19675.4]
  wire [7:0] _T_24993; // @[Mux.scala 19:72:@19682.4]
  wire [7:0] _T_25000; // @[Mux.scala 19:72:@19689.4]
  wire [15:0] _T_25001; // @[Mux.scala 19:72:@19690.4]
  wire [15:0] _T_25003; // @[Mux.scala 19:72:@19691.4]
  wire [15:0] _T_25018; // @[Mux.scala 19:72:@19706.4]
  wire [15:0] _T_25020; // @[Mux.scala 19:72:@19707.4]
  wire [15:0] _T_25035; // @[Mux.scala 19:72:@19722.4]
  wire [15:0] _T_25037; // @[Mux.scala 19:72:@19723.4]
  wire [15:0] _T_25052; // @[Mux.scala 19:72:@19738.4]
  wire [15:0] _T_25054; // @[Mux.scala 19:72:@19739.4]
  wire [15:0] _T_25069; // @[Mux.scala 19:72:@19754.4]
  wire [15:0] _T_25071; // @[Mux.scala 19:72:@19755.4]
  wire [15:0] _T_25086; // @[Mux.scala 19:72:@19770.4]
  wire [15:0] _T_25088; // @[Mux.scala 19:72:@19771.4]
  wire [15:0] _T_25103; // @[Mux.scala 19:72:@19786.4]
  wire [15:0] _T_25105; // @[Mux.scala 19:72:@19787.4]
  wire [15:0] _T_25120; // @[Mux.scala 19:72:@19802.4]
  wire [15:0] _T_25122; // @[Mux.scala 19:72:@19803.4]
  wire [15:0] _T_25137; // @[Mux.scala 19:72:@19818.4]
  wire [15:0] _T_25139; // @[Mux.scala 19:72:@19819.4]
  wire [15:0] _T_25140; // @[Mux.scala 19:72:@19820.4]
  wire [15:0] _T_25141; // @[Mux.scala 19:72:@19821.4]
  wire [15:0] _T_25142; // @[Mux.scala 19:72:@19822.4]
  wire [15:0] _T_25143; // @[Mux.scala 19:72:@19823.4]
  wire [15:0] _T_25144; // @[Mux.scala 19:72:@19824.4]
  wire [15:0] _T_25145; // @[Mux.scala 19:72:@19825.4]
  wire [15:0] _T_25146; // @[Mux.scala 19:72:@19826.4]
  wire [15:0] _T_25147; // @[Mux.scala 19:72:@19827.4]
  wire [15:0] _T_25148; // @[Mux.scala 19:72:@19828.4]
  wire [15:0] _T_25149; // @[Mux.scala 19:72:@19829.4]
  wire [15:0] _T_25150; // @[Mux.scala 19:72:@19830.4]
  wire [15:0] _T_25151; // @[Mux.scala 19:72:@19831.4]
  wire [15:0] _T_25152; // @[Mux.scala 19:72:@19832.4]
  wire [15:0] _T_25153; // @[Mux.scala 19:72:@19833.4]
  wire [15:0] _T_25154; // @[Mux.scala 19:72:@19834.4]
  wire [7:0] _T_25732; // @[Mux.scala 19:72:@20184.4]
  wire [7:0] _T_25739; // @[Mux.scala 19:72:@20191.4]
  wire [15:0] _T_25740; // @[Mux.scala 19:72:@20192.4]
  wire [15:0] _T_25742; // @[Mux.scala 19:72:@20193.4]
  wire [7:0] _T_25749; // @[Mux.scala 19:72:@20200.4]
  wire [7:0] _T_25756; // @[Mux.scala 19:72:@20207.4]
  wire [15:0] _T_25757; // @[Mux.scala 19:72:@20208.4]
  wire [15:0] _T_25759; // @[Mux.scala 19:72:@20209.4]
  wire [7:0] _T_25766; // @[Mux.scala 19:72:@20216.4]
  wire [7:0] _T_25773; // @[Mux.scala 19:72:@20223.4]
  wire [15:0] _T_25774; // @[Mux.scala 19:72:@20224.4]
  wire [15:0] _T_25776; // @[Mux.scala 19:72:@20225.4]
  wire [7:0] _T_25783; // @[Mux.scala 19:72:@20232.4]
  wire [7:0] _T_25790; // @[Mux.scala 19:72:@20239.4]
  wire [15:0] _T_25791; // @[Mux.scala 19:72:@20240.4]
  wire [15:0] _T_25793; // @[Mux.scala 19:72:@20241.4]
  wire [7:0] _T_25800; // @[Mux.scala 19:72:@20248.4]
  wire [7:0] _T_25807; // @[Mux.scala 19:72:@20255.4]
  wire [15:0] _T_25808; // @[Mux.scala 19:72:@20256.4]
  wire [15:0] _T_25810; // @[Mux.scala 19:72:@20257.4]
  wire [7:0] _T_25817; // @[Mux.scala 19:72:@20264.4]
  wire [7:0] _T_25824; // @[Mux.scala 19:72:@20271.4]
  wire [15:0] _T_25825; // @[Mux.scala 19:72:@20272.4]
  wire [15:0] _T_25827; // @[Mux.scala 19:72:@20273.4]
  wire [7:0] _T_25834; // @[Mux.scala 19:72:@20280.4]
  wire [7:0] _T_25841; // @[Mux.scala 19:72:@20287.4]
  wire [15:0] _T_25842; // @[Mux.scala 19:72:@20288.4]
  wire [15:0] _T_25844; // @[Mux.scala 19:72:@20289.4]
  wire [7:0] _T_25851; // @[Mux.scala 19:72:@20296.4]
  wire [7:0] _T_25858; // @[Mux.scala 19:72:@20303.4]
  wire [15:0] _T_25859; // @[Mux.scala 19:72:@20304.4]
  wire [15:0] _T_25861; // @[Mux.scala 19:72:@20305.4]
  wire [15:0] _T_25876; // @[Mux.scala 19:72:@20320.4]
  wire [15:0] _T_25878; // @[Mux.scala 19:72:@20321.4]
  wire [15:0] _T_25893; // @[Mux.scala 19:72:@20336.4]
  wire [15:0] _T_25895; // @[Mux.scala 19:72:@20337.4]
  wire [15:0] _T_25910; // @[Mux.scala 19:72:@20352.4]
  wire [15:0] _T_25912; // @[Mux.scala 19:72:@20353.4]
  wire [15:0] _T_25927; // @[Mux.scala 19:72:@20368.4]
  wire [15:0] _T_25929; // @[Mux.scala 19:72:@20369.4]
  wire [15:0] _T_25944; // @[Mux.scala 19:72:@20384.4]
  wire [15:0] _T_25946; // @[Mux.scala 19:72:@20385.4]
  wire [15:0] _T_25961; // @[Mux.scala 19:72:@20400.4]
  wire [15:0] _T_25963; // @[Mux.scala 19:72:@20401.4]
  wire [15:0] _T_25978; // @[Mux.scala 19:72:@20416.4]
  wire [15:0] _T_25980; // @[Mux.scala 19:72:@20417.4]
  wire [15:0] _T_25995; // @[Mux.scala 19:72:@20432.4]
  wire [15:0] _T_25997; // @[Mux.scala 19:72:@20433.4]
  wire [15:0] _T_25998; // @[Mux.scala 19:72:@20434.4]
  wire [15:0] _T_25999; // @[Mux.scala 19:72:@20435.4]
  wire [15:0] _T_26000; // @[Mux.scala 19:72:@20436.4]
  wire [15:0] _T_26001; // @[Mux.scala 19:72:@20437.4]
  wire [15:0] _T_26002; // @[Mux.scala 19:72:@20438.4]
  wire [15:0] _T_26003; // @[Mux.scala 19:72:@20439.4]
  wire [15:0] _T_26004; // @[Mux.scala 19:72:@20440.4]
  wire [15:0] _T_26005; // @[Mux.scala 19:72:@20441.4]
  wire [15:0] _T_26006; // @[Mux.scala 19:72:@20442.4]
  wire [15:0] _T_26007; // @[Mux.scala 19:72:@20443.4]
  wire [15:0] _T_26008; // @[Mux.scala 19:72:@20444.4]
  wire [15:0] _T_26009; // @[Mux.scala 19:72:@20445.4]
  wire [15:0] _T_26010; // @[Mux.scala 19:72:@20446.4]
  wire [15:0] _T_26011; // @[Mux.scala 19:72:@20447.4]
  wire [15:0] _T_26012; // @[Mux.scala 19:72:@20448.4]
  wire [7:0] _T_26590; // @[Mux.scala 19:72:@20798.4]
  wire [7:0] _T_26597; // @[Mux.scala 19:72:@20805.4]
  wire [15:0] _T_26598; // @[Mux.scala 19:72:@20806.4]
  wire [15:0] _T_26600; // @[Mux.scala 19:72:@20807.4]
  wire [7:0] _T_26607; // @[Mux.scala 19:72:@20814.4]
  wire [7:0] _T_26614; // @[Mux.scala 19:72:@20821.4]
  wire [15:0] _T_26615; // @[Mux.scala 19:72:@20822.4]
  wire [15:0] _T_26617; // @[Mux.scala 19:72:@20823.4]
  wire [7:0] _T_26624; // @[Mux.scala 19:72:@20830.4]
  wire [7:0] _T_26631; // @[Mux.scala 19:72:@20837.4]
  wire [15:0] _T_26632; // @[Mux.scala 19:72:@20838.4]
  wire [15:0] _T_26634; // @[Mux.scala 19:72:@20839.4]
  wire [7:0] _T_26641; // @[Mux.scala 19:72:@20846.4]
  wire [7:0] _T_26648; // @[Mux.scala 19:72:@20853.4]
  wire [15:0] _T_26649; // @[Mux.scala 19:72:@20854.4]
  wire [15:0] _T_26651; // @[Mux.scala 19:72:@20855.4]
  wire [7:0] _T_26658; // @[Mux.scala 19:72:@20862.4]
  wire [7:0] _T_26665; // @[Mux.scala 19:72:@20869.4]
  wire [15:0] _T_26666; // @[Mux.scala 19:72:@20870.4]
  wire [15:0] _T_26668; // @[Mux.scala 19:72:@20871.4]
  wire [7:0] _T_26675; // @[Mux.scala 19:72:@20878.4]
  wire [7:0] _T_26682; // @[Mux.scala 19:72:@20885.4]
  wire [15:0] _T_26683; // @[Mux.scala 19:72:@20886.4]
  wire [15:0] _T_26685; // @[Mux.scala 19:72:@20887.4]
  wire [7:0] _T_26692; // @[Mux.scala 19:72:@20894.4]
  wire [7:0] _T_26699; // @[Mux.scala 19:72:@20901.4]
  wire [15:0] _T_26700; // @[Mux.scala 19:72:@20902.4]
  wire [15:0] _T_26702; // @[Mux.scala 19:72:@20903.4]
  wire [7:0] _T_26709; // @[Mux.scala 19:72:@20910.4]
  wire [7:0] _T_26716; // @[Mux.scala 19:72:@20917.4]
  wire [15:0] _T_26717; // @[Mux.scala 19:72:@20918.4]
  wire [15:0] _T_26719; // @[Mux.scala 19:72:@20919.4]
  wire [15:0] _T_26734; // @[Mux.scala 19:72:@20934.4]
  wire [15:0] _T_26736; // @[Mux.scala 19:72:@20935.4]
  wire [15:0] _T_26751; // @[Mux.scala 19:72:@20950.4]
  wire [15:0] _T_26753; // @[Mux.scala 19:72:@20951.4]
  wire [15:0] _T_26768; // @[Mux.scala 19:72:@20966.4]
  wire [15:0] _T_26770; // @[Mux.scala 19:72:@20967.4]
  wire [15:0] _T_26785; // @[Mux.scala 19:72:@20982.4]
  wire [15:0] _T_26787; // @[Mux.scala 19:72:@20983.4]
  wire [15:0] _T_26802; // @[Mux.scala 19:72:@20998.4]
  wire [15:0] _T_26804; // @[Mux.scala 19:72:@20999.4]
  wire [15:0] _T_26819; // @[Mux.scala 19:72:@21014.4]
  wire [15:0] _T_26821; // @[Mux.scala 19:72:@21015.4]
  wire [15:0] _T_26836; // @[Mux.scala 19:72:@21030.4]
  wire [15:0] _T_26838; // @[Mux.scala 19:72:@21031.4]
  wire [15:0] _T_26853; // @[Mux.scala 19:72:@21046.4]
  wire [15:0] _T_26855; // @[Mux.scala 19:72:@21047.4]
  wire [15:0] _T_26856; // @[Mux.scala 19:72:@21048.4]
  wire [15:0] _T_26857; // @[Mux.scala 19:72:@21049.4]
  wire [15:0] _T_26858; // @[Mux.scala 19:72:@21050.4]
  wire [15:0] _T_26859; // @[Mux.scala 19:72:@21051.4]
  wire [15:0] _T_26860; // @[Mux.scala 19:72:@21052.4]
  wire [15:0] _T_26861; // @[Mux.scala 19:72:@21053.4]
  wire [15:0] _T_26862; // @[Mux.scala 19:72:@21054.4]
  wire [15:0] _T_26863; // @[Mux.scala 19:72:@21055.4]
  wire [15:0] _T_26864; // @[Mux.scala 19:72:@21056.4]
  wire [15:0] _T_26865; // @[Mux.scala 19:72:@21057.4]
  wire [15:0] _T_26866; // @[Mux.scala 19:72:@21058.4]
  wire [15:0] _T_26867; // @[Mux.scala 19:72:@21059.4]
  wire [15:0] _T_26868; // @[Mux.scala 19:72:@21060.4]
  wire [15:0] _T_26869; // @[Mux.scala 19:72:@21061.4]
  wire [15:0] _T_26870; // @[Mux.scala 19:72:@21062.4]
  wire [7:0] _T_27448; // @[Mux.scala 19:72:@21412.4]
  wire [7:0] _T_27455; // @[Mux.scala 19:72:@21419.4]
  wire [15:0] _T_27456; // @[Mux.scala 19:72:@21420.4]
  wire [15:0] _T_27458; // @[Mux.scala 19:72:@21421.4]
  wire [7:0] _T_27465; // @[Mux.scala 19:72:@21428.4]
  wire [7:0] _T_27472; // @[Mux.scala 19:72:@21435.4]
  wire [15:0] _T_27473; // @[Mux.scala 19:72:@21436.4]
  wire [15:0] _T_27475; // @[Mux.scala 19:72:@21437.4]
  wire [7:0] _T_27482; // @[Mux.scala 19:72:@21444.4]
  wire [7:0] _T_27489; // @[Mux.scala 19:72:@21451.4]
  wire [15:0] _T_27490; // @[Mux.scala 19:72:@21452.4]
  wire [15:0] _T_27492; // @[Mux.scala 19:72:@21453.4]
  wire [7:0] _T_27499; // @[Mux.scala 19:72:@21460.4]
  wire [7:0] _T_27506; // @[Mux.scala 19:72:@21467.4]
  wire [15:0] _T_27507; // @[Mux.scala 19:72:@21468.4]
  wire [15:0] _T_27509; // @[Mux.scala 19:72:@21469.4]
  wire [7:0] _T_27516; // @[Mux.scala 19:72:@21476.4]
  wire [7:0] _T_27523; // @[Mux.scala 19:72:@21483.4]
  wire [15:0] _T_27524; // @[Mux.scala 19:72:@21484.4]
  wire [15:0] _T_27526; // @[Mux.scala 19:72:@21485.4]
  wire [7:0] _T_27533; // @[Mux.scala 19:72:@21492.4]
  wire [7:0] _T_27540; // @[Mux.scala 19:72:@21499.4]
  wire [15:0] _T_27541; // @[Mux.scala 19:72:@21500.4]
  wire [15:0] _T_27543; // @[Mux.scala 19:72:@21501.4]
  wire [7:0] _T_27550; // @[Mux.scala 19:72:@21508.4]
  wire [7:0] _T_27557; // @[Mux.scala 19:72:@21515.4]
  wire [15:0] _T_27558; // @[Mux.scala 19:72:@21516.4]
  wire [15:0] _T_27560; // @[Mux.scala 19:72:@21517.4]
  wire [7:0] _T_27567; // @[Mux.scala 19:72:@21524.4]
  wire [7:0] _T_27574; // @[Mux.scala 19:72:@21531.4]
  wire [15:0] _T_27575; // @[Mux.scala 19:72:@21532.4]
  wire [15:0] _T_27577; // @[Mux.scala 19:72:@21533.4]
  wire [15:0] _T_27592; // @[Mux.scala 19:72:@21548.4]
  wire [15:0] _T_27594; // @[Mux.scala 19:72:@21549.4]
  wire [15:0] _T_27609; // @[Mux.scala 19:72:@21564.4]
  wire [15:0] _T_27611; // @[Mux.scala 19:72:@21565.4]
  wire [15:0] _T_27626; // @[Mux.scala 19:72:@21580.4]
  wire [15:0] _T_27628; // @[Mux.scala 19:72:@21581.4]
  wire [15:0] _T_27643; // @[Mux.scala 19:72:@21596.4]
  wire [15:0] _T_27645; // @[Mux.scala 19:72:@21597.4]
  wire [15:0] _T_27660; // @[Mux.scala 19:72:@21612.4]
  wire [15:0] _T_27662; // @[Mux.scala 19:72:@21613.4]
  wire [15:0] _T_27677; // @[Mux.scala 19:72:@21628.4]
  wire [15:0] _T_27679; // @[Mux.scala 19:72:@21629.4]
  wire [15:0] _T_27694; // @[Mux.scala 19:72:@21644.4]
  wire [15:0] _T_27696; // @[Mux.scala 19:72:@21645.4]
  wire [15:0] _T_27711; // @[Mux.scala 19:72:@21660.4]
  wire [15:0] _T_27713; // @[Mux.scala 19:72:@21661.4]
  wire [15:0] _T_27714; // @[Mux.scala 19:72:@21662.4]
  wire [15:0] _T_27715; // @[Mux.scala 19:72:@21663.4]
  wire [15:0] _T_27716; // @[Mux.scala 19:72:@21664.4]
  wire [15:0] _T_27717; // @[Mux.scala 19:72:@21665.4]
  wire [15:0] _T_27718; // @[Mux.scala 19:72:@21666.4]
  wire [15:0] _T_27719; // @[Mux.scala 19:72:@21667.4]
  wire [15:0] _T_27720; // @[Mux.scala 19:72:@21668.4]
  wire [15:0] _T_27721; // @[Mux.scala 19:72:@21669.4]
  wire [15:0] _T_27722; // @[Mux.scala 19:72:@21670.4]
  wire [15:0] _T_27723; // @[Mux.scala 19:72:@21671.4]
  wire [15:0] _T_27724; // @[Mux.scala 19:72:@21672.4]
  wire [15:0] _T_27725; // @[Mux.scala 19:72:@21673.4]
  wire [15:0] _T_27726; // @[Mux.scala 19:72:@21674.4]
  wire [15:0] _T_27727; // @[Mux.scala 19:72:@21675.4]
  wire [15:0] _T_27728; // @[Mux.scala 19:72:@21676.4]
  wire [7:0] _T_28306; // @[Mux.scala 19:72:@22026.4]
  wire [7:0] _T_28313; // @[Mux.scala 19:72:@22033.4]
  wire [15:0] _T_28314; // @[Mux.scala 19:72:@22034.4]
  wire [15:0] _T_28316; // @[Mux.scala 19:72:@22035.4]
  wire [7:0] _T_28323; // @[Mux.scala 19:72:@22042.4]
  wire [7:0] _T_28330; // @[Mux.scala 19:72:@22049.4]
  wire [15:0] _T_28331; // @[Mux.scala 19:72:@22050.4]
  wire [15:0] _T_28333; // @[Mux.scala 19:72:@22051.4]
  wire [7:0] _T_28340; // @[Mux.scala 19:72:@22058.4]
  wire [7:0] _T_28347; // @[Mux.scala 19:72:@22065.4]
  wire [15:0] _T_28348; // @[Mux.scala 19:72:@22066.4]
  wire [15:0] _T_28350; // @[Mux.scala 19:72:@22067.4]
  wire [7:0] _T_28357; // @[Mux.scala 19:72:@22074.4]
  wire [7:0] _T_28364; // @[Mux.scala 19:72:@22081.4]
  wire [15:0] _T_28365; // @[Mux.scala 19:72:@22082.4]
  wire [15:0] _T_28367; // @[Mux.scala 19:72:@22083.4]
  wire [7:0] _T_28374; // @[Mux.scala 19:72:@22090.4]
  wire [7:0] _T_28381; // @[Mux.scala 19:72:@22097.4]
  wire [15:0] _T_28382; // @[Mux.scala 19:72:@22098.4]
  wire [15:0] _T_28384; // @[Mux.scala 19:72:@22099.4]
  wire [7:0] _T_28391; // @[Mux.scala 19:72:@22106.4]
  wire [7:0] _T_28398; // @[Mux.scala 19:72:@22113.4]
  wire [15:0] _T_28399; // @[Mux.scala 19:72:@22114.4]
  wire [15:0] _T_28401; // @[Mux.scala 19:72:@22115.4]
  wire [7:0] _T_28408; // @[Mux.scala 19:72:@22122.4]
  wire [7:0] _T_28415; // @[Mux.scala 19:72:@22129.4]
  wire [15:0] _T_28416; // @[Mux.scala 19:72:@22130.4]
  wire [15:0] _T_28418; // @[Mux.scala 19:72:@22131.4]
  wire [7:0] _T_28425; // @[Mux.scala 19:72:@22138.4]
  wire [7:0] _T_28432; // @[Mux.scala 19:72:@22145.4]
  wire [15:0] _T_28433; // @[Mux.scala 19:72:@22146.4]
  wire [15:0] _T_28435; // @[Mux.scala 19:72:@22147.4]
  wire [15:0] _T_28450; // @[Mux.scala 19:72:@22162.4]
  wire [15:0] _T_28452; // @[Mux.scala 19:72:@22163.4]
  wire [15:0] _T_28467; // @[Mux.scala 19:72:@22178.4]
  wire [15:0] _T_28469; // @[Mux.scala 19:72:@22179.4]
  wire [15:0] _T_28484; // @[Mux.scala 19:72:@22194.4]
  wire [15:0] _T_28486; // @[Mux.scala 19:72:@22195.4]
  wire [15:0] _T_28501; // @[Mux.scala 19:72:@22210.4]
  wire [15:0] _T_28503; // @[Mux.scala 19:72:@22211.4]
  wire [15:0] _T_28518; // @[Mux.scala 19:72:@22226.4]
  wire [15:0] _T_28520; // @[Mux.scala 19:72:@22227.4]
  wire [15:0] _T_28535; // @[Mux.scala 19:72:@22242.4]
  wire [15:0] _T_28537; // @[Mux.scala 19:72:@22243.4]
  wire [15:0] _T_28552; // @[Mux.scala 19:72:@22258.4]
  wire [15:0] _T_28554; // @[Mux.scala 19:72:@22259.4]
  wire [15:0] _T_28569; // @[Mux.scala 19:72:@22274.4]
  wire [15:0] _T_28571; // @[Mux.scala 19:72:@22275.4]
  wire [15:0] _T_28572; // @[Mux.scala 19:72:@22276.4]
  wire [15:0] _T_28573; // @[Mux.scala 19:72:@22277.4]
  wire [15:0] _T_28574; // @[Mux.scala 19:72:@22278.4]
  wire [15:0] _T_28575; // @[Mux.scala 19:72:@22279.4]
  wire [15:0] _T_28576; // @[Mux.scala 19:72:@22280.4]
  wire [15:0] _T_28577; // @[Mux.scala 19:72:@22281.4]
  wire [15:0] _T_28578; // @[Mux.scala 19:72:@22282.4]
  wire [15:0] _T_28579; // @[Mux.scala 19:72:@22283.4]
  wire [15:0] _T_28580; // @[Mux.scala 19:72:@22284.4]
  wire [15:0] _T_28581; // @[Mux.scala 19:72:@22285.4]
  wire [15:0] _T_28582; // @[Mux.scala 19:72:@22286.4]
  wire [15:0] _T_28583; // @[Mux.scala 19:72:@22287.4]
  wire [15:0] _T_28584; // @[Mux.scala 19:72:@22288.4]
  wire [15:0] _T_28585; // @[Mux.scala 19:72:@22289.4]
  wire [15:0] _T_28586; // @[Mux.scala 19:72:@22290.4]
  wire [7:0] _T_29164; // @[Mux.scala 19:72:@22640.4]
  wire [7:0] _T_29171; // @[Mux.scala 19:72:@22647.4]
  wire [15:0] _T_29172; // @[Mux.scala 19:72:@22648.4]
  wire [15:0] _T_29174; // @[Mux.scala 19:72:@22649.4]
  wire [7:0] _T_29181; // @[Mux.scala 19:72:@22656.4]
  wire [7:0] _T_29188; // @[Mux.scala 19:72:@22663.4]
  wire [15:0] _T_29189; // @[Mux.scala 19:72:@22664.4]
  wire [15:0] _T_29191; // @[Mux.scala 19:72:@22665.4]
  wire [7:0] _T_29198; // @[Mux.scala 19:72:@22672.4]
  wire [7:0] _T_29205; // @[Mux.scala 19:72:@22679.4]
  wire [15:0] _T_29206; // @[Mux.scala 19:72:@22680.4]
  wire [15:0] _T_29208; // @[Mux.scala 19:72:@22681.4]
  wire [7:0] _T_29215; // @[Mux.scala 19:72:@22688.4]
  wire [7:0] _T_29222; // @[Mux.scala 19:72:@22695.4]
  wire [15:0] _T_29223; // @[Mux.scala 19:72:@22696.4]
  wire [15:0] _T_29225; // @[Mux.scala 19:72:@22697.4]
  wire [7:0] _T_29232; // @[Mux.scala 19:72:@22704.4]
  wire [7:0] _T_29239; // @[Mux.scala 19:72:@22711.4]
  wire [15:0] _T_29240; // @[Mux.scala 19:72:@22712.4]
  wire [15:0] _T_29242; // @[Mux.scala 19:72:@22713.4]
  wire [7:0] _T_29249; // @[Mux.scala 19:72:@22720.4]
  wire [7:0] _T_29256; // @[Mux.scala 19:72:@22727.4]
  wire [15:0] _T_29257; // @[Mux.scala 19:72:@22728.4]
  wire [15:0] _T_29259; // @[Mux.scala 19:72:@22729.4]
  wire [7:0] _T_29266; // @[Mux.scala 19:72:@22736.4]
  wire [7:0] _T_29273; // @[Mux.scala 19:72:@22743.4]
  wire [15:0] _T_29274; // @[Mux.scala 19:72:@22744.4]
  wire [15:0] _T_29276; // @[Mux.scala 19:72:@22745.4]
  wire [7:0] _T_29283; // @[Mux.scala 19:72:@22752.4]
  wire [7:0] _T_29290; // @[Mux.scala 19:72:@22759.4]
  wire [15:0] _T_29291; // @[Mux.scala 19:72:@22760.4]
  wire [15:0] _T_29293; // @[Mux.scala 19:72:@22761.4]
  wire [15:0] _T_29308; // @[Mux.scala 19:72:@22776.4]
  wire [15:0] _T_29310; // @[Mux.scala 19:72:@22777.4]
  wire [15:0] _T_29325; // @[Mux.scala 19:72:@22792.4]
  wire [15:0] _T_29327; // @[Mux.scala 19:72:@22793.4]
  wire [15:0] _T_29342; // @[Mux.scala 19:72:@22808.4]
  wire [15:0] _T_29344; // @[Mux.scala 19:72:@22809.4]
  wire [15:0] _T_29359; // @[Mux.scala 19:72:@22824.4]
  wire [15:0] _T_29361; // @[Mux.scala 19:72:@22825.4]
  wire [15:0] _T_29376; // @[Mux.scala 19:72:@22840.4]
  wire [15:0] _T_29378; // @[Mux.scala 19:72:@22841.4]
  wire [15:0] _T_29393; // @[Mux.scala 19:72:@22856.4]
  wire [15:0] _T_29395; // @[Mux.scala 19:72:@22857.4]
  wire [15:0] _T_29410; // @[Mux.scala 19:72:@22872.4]
  wire [15:0] _T_29412; // @[Mux.scala 19:72:@22873.4]
  wire [15:0] _T_29427; // @[Mux.scala 19:72:@22888.4]
  wire [15:0] _T_29429; // @[Mux.scala 19:72:@22889.4]
  wire [15:0] _T_29430; // @[Mux.scala 19:72:@22890.4]
  wire [15:0] _T_29431; // @[Mux.scala 19:72:@22891.4]
  wire [15:0] _T_29432; // @[Mux.scala 19:72:@22892.4]
  wire [15:0] _T_29433; // @[Mux.scala 19:72:@22893.4]
  wire [15:0] _T_29434; // @[Mux.scala 19:72:@22894.4]
  wire [15:0] _T_29435; // @[Mux.scala 19:72:@22895.4]
  wire [15:0] _T_29436; // @[Mux.scala 19:72:@22896.4]
  wire [15:0] _T_29437; // @[Mux.scala 19:72:@22897.4]
  wire [15:0] _T_29438; // @[Mux.scala 19:72:@22898.4]
  wire [15:0] _T_29439; // @[Mux.scala 19:72:@22899.4]
  wire [15:0] _T_29440; // @[Mux.scala 19:72:@22900.4]
  wire [15:0] _T_29441; // @[Mux.scala 19:72:@22901.4]
  wire [15:0] _T_29442; // @[Mux.scala 19:72:@22902.4]
  wire [15:0] _T_29443; // @[Mux.scala 19:72:@22903.4]
  wire [15:0] _T_29444; // @[Mux.scala 19:72:@22904.4]
  wire [7:0] _T_30022; // @[Mux.scala 19:72:@23254.4]
  wire [7:0] _T_30029; // @[Mux.scala 19:72:@23261.4]
  wire [15:0] _T_30030; // @[Mux.scala 19:72:@23262.4]
  wire [15:0] _T_30032; // @[Mux.scala 19:72:@23263.4]
  wire [7:0] _T_30039; // @[Mux.scala 19:72:@23270.4]
  wire [7:0] _T_30046; // @[Mux.scala 19:72:@23277.4]
  wire [15:0] _T_30047; // @[Mux.scala 19:72:@23278.4]
  wire [15:0] _T_30049; // @[Mux.scala 19:72:@23279.4]
  wire [7:0] _T_30056; // @[Mux.scala 19:72:@23286.4]
  wire [7:0] _T_30063; // @[Mux.scala 19:72:@23293.4]
  wire [15:0] _T_30064; // @[Mux.scala 19:72:@23294.4]
  wire [15:0] _T_30066; // @[Mux.scala 19:72:@23295.4]
  wire [7:0] _T_30073; // @[Mux.scala 19:72:@23302.4]
  wire [7:0] _T_30080; // @[Mux.scala 19:72:@23309.4]
  wire [15:0] _T_30081; // @[Mux.scala 19:72:@23310.4]
  wire [15:0] _T_30083; // @[Mux.scala 19:72:@23311.4]
  wire [7:0] _T_30090; // @[Mux.scala 19:72:@23318.4]
  wire [7:0] _T_30097; // @[Mux.scala 19:72:@23325.4]
  wire [15:0] _T_30098; // @[Mux.scala 19:72:@23326.4]
  wire [15:0] _T_30100; // @[Mux.scala 19:72:@23327.4]
  wire [7:0] _T_30107; // @[Mux.scala 19:72:@23334.4]
  wire [7:0] _T_30114; // @[Mux.scala 19:72:@23341.4]
  wire [15:0] _T_30115; // @[Mux.scala 19:72:@23342.4]
  wire [15:0] _T_30117; // @[Mux.scala 19:72:@23343.4]
  wire [7:0] _T_30124; // @[Mux.scala 19:72:@23350.4]
  wire [7:0] _T_30131; // @[Mux.scala 19:72:@23357.4]
  wire [15:0] _T_30132; // @[Mux.scala 19:72:@23358.4]
  wire [15:0] _T_30134; // @[Mux.scala 19:72:@23359.4]
  wire [7:0] _T_30141; // @[Mux.scala 19:72:@23366.4]
  wire [7:0] _T_30148; // @[Mux.scala 19:72:@23373.4]
  wire [15:0] _T_30149; // @[Mux.scala 19:72:@23374.4]
  wire [15:0] _T_30151; // @[Mux.scala 19:72:@23375.4]
  wire [15:0] _T_30166; // @[Mux.scala 19:72:@23390.4]
  wire [15:0] _T_30168; // @[Mux.scala 19:72:@23391.4]
  wire [15:0] _T_30183; // @[Mux.scala 19:72:@23406.4]
  wire [15:0] _T_30185; // @[Mux.scala 19:72:@23407.4]
  wire [15:0] _T_30200; // @[Mux.scala 19:72:@23422.4]
  wire [15:0] _T_30202; // @[Mux.scala 19:72:@23423.4]
  wire [15:0] _T_30217; // @[Mux.scala 19:72:@23438.4]
  wire [15:0] _T_30219; // @[Mux.scala 19:72:@23439.4]
  wire [15:0] _T_30234; // @[Mux.scala 19:72:@23454.4]
  wire [15:0] _T_30236; // @[Mux.scala 19:72:@23455.4]
  wire [15:0] _T_30251; // @[Mux.scala 19:72:@23470.4]
  wire [15:0] _T_30253; // @[Mux.scala 19:72:@23471.4]
  wire [15:0] _T_30268; // @[Mux.scala 19:72:@23486.4]
  wire [15:0] _T_30270; // @[Mux.scala 19:72:@23487.4]
  wire [15:0] _T_30285; // @[Mux.scala 19:72:@23502.4]
  wire [15:0] _T_30287; // @[Mux.scala 19:72:@23503.4]
  wire [15:0] _T_30288; // @[Mux.scala 19:72:@23504.4]
  wire [15:0] _T_30289; // @[Mux.scala 19:72:@23505.4]
  wire [15:0] _T_30290; // @[Mux.scala 19:72:@23506.4]
  wire [15:0] _T_30291; // @[Mux.scala 19:72:@23507.4]
  wire [15:0] _T_30292; // @[Mux.scala 19:72:@23508.4]
  wire [15:0] _T_30293; // @[Mux.scala 19:72:@23509.4]
  wire [15:0] _T_30294; // @[Mux.scala 19:72:@23510.4]
  wire [15:0] _T_30295; // @[Mux.scala 19:72:@23511.4]
  wire [15:0] _T_30296; // @[Mux.scala 19:72:@23512.4]
  wire [15:0] _T_30297; // @[Mux.scala 19:72:@23513.4]
  wire [15:0] _T_30298; // @[Mux.scala 19:72:@23514.4]
  wire [15:0] _T_30299; // @[Mux.scala 19:72:@23515.4]
  wire [15:0] _T_30300; // @[Mux.scala 19:72:@23516.4]
  wire [15:0] _T_30301; // @[Mux.scala 19:72:@23517.4]
  wire [15:0] _T_30302; // @[Mux.scala 19:72:@23518.4]
  wire [7:0] _T_30880; // @[Mux.scala 19:72:@23868.4]
  wire [7:0] _T_30887; // @[Mux.scala 19:72:@23875.4]
  wire [15:0] _T_30888; // @[Mux.scala 19:72:@23876.4]
  wire [15:0] _T_30890; // @[Mux.scala 19:72:@23877.4]
  wire [7:0] _T_30897; // @[Mux.scala 19:72:@23884.4]
  wire [7:0] _T_30904; // @[Mux.scala 19:72:@23891.4]
  wire [15:0] _T_30905; // @[Mux.scala 19:72:@23892.4]
  wire [15:0] _T_30907; // @[Mux.scala 19:72:@23893.4]
  wire [7:0] _T_30914; // @[Mux.scala 19:72:@23900.4]
  wire [7:0] _T_30921; // @[Mux.scala 19:72:@23907.4]
  wire [15:0] _T_30922; // @[Mux.scala 19:72:@23908.4]
  wire [15:0] _T_30924; // @[Mux.scala 19:72:@23909.4]
  wire [7:0] _T_30931; // @[Mux.scala 19:72:@23916.4]
  wire [7:0] _T_30938; // @[Mux.scala 19:72:@23923.4]
  wire [15:0] _T_30939; // @[Mux.scala 19:72:@23924.4]
  wire [15:0] _T_30941; // @[Mux.scala 19:72:@23925.4]
  wire [7:0] _T_30948; // @[Mux.scala 19:72:@23932.4]
  wire [7:0] _T_30955; // @[Mux.scala 19:72:@23939.4]
  wire [15:0] _T_30956; // @[Mux.scala 19:72:@23940.4]
  wire [15:0] _T_30958; // @[Mux.scala 19:72:@23941.4]
  wire [7:0] _T_30965; // @[Mux.scala 19:72:@23948.4]
  wire [7:0] _T_30972; // @[Mux.scala 19:72:@23955.4]
  wire [15:0] _T_30973; // @[Mux.scala 19:72:@23956.4]
  wire [15:0] _T_30975; // @[Mux.scala 19:72:@23957.4]
  wire [7:0] _T_30982; // @[Mux.scala 19:72:@23964.4]
  wire [7:0] _T_30989; // @[Mux.scala 19:72:@23971.4]
  wire [15:0] _T_30990; // @[Mux.scala 19:72:@23972.4]
  wire [15:0] _T_30992; // @[Mux.scala 19:72:@23973.4]
  wire [7:0] _T_30999; // @[Mux.scala 19:72:@23980.4]
  wire [7:0] _T_31006; // @[Mux.scala 19:72:@23987.4]
  wire [15:0] _T_31007; // @[Mux.scala 19:72:@23988.4]
  wire [15:0] _T_31009; // @[Mux.scala 19:72:@23989.4]
  wire [15:0] _T_31024; // @[Mux.scala 19:72:@24004.4]
  wire [15:0] _T_31026; // @[Mux.scala 19:72:@24005.4]
  wire [15:0] _T_31041; // @[Mux.scala 19:72:@24020.4]
  wire [15:0] _T_31043; // @[Mux.scala 19:72:@24021.4]
  wire [15:0] _T_31058; // @[Mux.scala 19:72:@24036.4]
  wire [15:0] _T_31060; // @[Mux.scala 19:72:@24037.4]
  wire [15:0] _T_31075; // @[Mux.scala 19:72:@24052.4]
  wire [15:0] _T_31077; // @[Mux.scala 19:72:@24053.4]
  wire [15:0] _T_31092; // @[Mux.scala 19:72:@24068.4]
  wire [15:0] _T_31094; // @[Mux.scala 19:72:@24069.4]
  wire [15:0] _T_31109; // @[Mux.scala 19:72:@24084.4]
  wire [15:0] _T_31111; // @[Mux.scala 19:72:@24085.4]
  wire [15:0] _T_31126; // @[Mux.scala 19:72:@24100.4]
  wire [15:0] _T_31128; // @[Mux.scala 19:72:@24101.4]
  wire [15:0] _T_31143; // @[Mux.scala 19:72:@24116.4]
  wire [15:0] _T_31145; // @[Mux.scala 19:72:@24117.4]
  wire [15:0] _T_31146; // @[Mux.scala 19:72:@24118.4]
  wire [15:0] _T_31147; // @[Mux.scala 19:72:@24119.4]
  wire [15:0] _T_31148; // @[Mux.scala 19:72:@24120.4]
  wire [15:0] _T_31149; // @[Mux.scala 19:72:@24121.4]
  wire [15:0] _T_31150; // @[Mux.scala 19:72:@24122.4]
  wire [15:0] _T_31151; // @[Mux.scala 19:72:@24123.4]
  wire [15:0] _T_31152; // @[Mux.scala 19:72:@24124.4]
  wire [15:0] _T_31153; // @[Mux.scala 19:72:@24125.4]
  wire [15:0] _T_31154; // @[Mux.scala 19:72:@24126.4]
  wire [15:0] _T_31155; // @[Mux.scala 19:72:@24127.4]
  wire [15:0] _T_31156; // @[Mux.scala 19:72:@24128.4]
  wire [15:0] _T_31157; // @[Mux.scala 19:72:@24129.4]
  wire [15:0] _T_31158; // @[Mux.scala 19:72:@24130.4]
  wire [15:0] _T_31159; // @[Mux.scala 19:72:@24131.4]
  wire [15:0] _T_31160; // @[Mux.scala 19:72:@24132.4]
  reg  conflictPReg_0_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_163;
  reg  conflictPReg_0_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_164;
  reg  conflictPReg_0_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_165;
  reg  conflictPReg_0_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_166;
  reg  conflictPReg_0_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_167;
  reg  conflictPReg_0_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_168;
  reg  conflictPReg_0_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_169;
  reg  conflictPReg_0_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_170;
  reg  conflictPReg_0_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_171;
  reg  conflictPReg_0_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_172;
  reg  conflictPReg_0_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_173;
  reg  conflictPReg_0_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_174;
  reg  conflictPReg_0_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_175;
  reg  conflictPReg_0_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_176;
  reg  conflictPReg_0_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_177;
  reg  conflictPReg_0_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_178;
  reg  conflictPReg_1_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_179;
  reg  conflictPReg_1_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_180;
  reg  conflictPReg_1_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_181;
  reg  conflictPReg_1_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_182;
  reg  conflictPReg_1_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_183;
  reg  conflictPReg_1_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_184;
  reg  conflictPReg_1_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_185;
  reg  conflictPReg_1_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_186;
  reg  conflictPReg_1_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_187;
  reg  conflictPReg_1_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_188;
  reg  conflictPReg_1_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_189;
  reg  conflictPReg_1_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_190;
  reg  conflictPReg_1_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_191;
  reg  conflictPReg_1_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_192;
  reg  conflictPReg_1_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_193;
  reg  conflictPReg_1_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_194;
  reg  conflictPReg_2_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_195;
  reg  conflictPReg_2_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_196;
  reg  conflictPReg_2_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_197;
  reg  conflictPReg_2_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_198;
  reg  conflictPReg_2_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_199;
  reg  conflictPReg_2_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_200;
  reg  conflictPReg_2_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_201;
  reg  conflictPReg_2_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_202;
  reg  conflictPReg_2_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_203;
  reg  conflictPReg_2_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_204;
  reg  conflictPReg_2_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_205;
  reg  conflictPReg_2_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_206;
  reg  conflictPReg_2_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_207;
  reg  conflictPReg_2_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_208;
  reg  conflictPReg_2_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_209;
  reg  conflictPReg_2_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_210;
  reg  conflictPReg_3_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_211;
  reg  conflictPReg_3_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_212;
  reg  conflictPReg_3_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_213;
  reg  conflictPReg_3_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_214;
  reg  conflictPReg_3_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_215;
  reg  conflictPReg_3_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_216;
  reg  conflictPReg_3_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_217;
  reg  conflictPReg_3_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_218;
  reg  conflictPReg_3_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_219;
  reg  conflictPReg_3_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_220;
  reg  conflictPReg_3_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_221;
  reg  conflictPReg_3_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_222;
  reg  conflictPReg_3_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_223;
  reg  conflictPReg_3_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_224;
  reg  conflictPReg_3_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_225;
  reg  conflictPReg_3_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_226;
  reg  conflictPReg_4_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_227;
  reg  conflictPReg_4_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_228;
  reg  conflictPReg_4_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_229;
  reg  conflictPReg_4_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_230;
  reg  conflictPReg_4_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_231;
  reg  conflictPReg_4_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_232;
  reg  conflictPReg_4_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_233;
  reg  conflictPReg_4_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_234;
  reg  conflictPReg_4_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_235;
  reg  conflictPReg_4_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_236;
  reg  conflictPReg_4_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_237;
  reg  conflictPReg_4_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_238;
  reg  conflictPReg_4_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_239;
  reg  conflictPReg_4_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_240;
  reg  conflictPReg_4_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_241;
  reg  conflictPReg_4_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_242;
  reg  conflictPReg_5_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_243;
  reg  conflictPReg_5_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_244;
  reg  conflictPReg_5_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_245;
  reg  conflictPReg_5_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_246;
  reg  conflictPReg_5_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_247;
  reg  conflictPReg_5_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_248;
  reg  conflictPReg_5_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_249;
  reg  conflictPReg_5_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_250;
  reg  conflictPReg_5_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_251;
  reg  conflictPReg_5_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_252;
  reg  conflictPReg_5_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_253;
  reg  conflictPReg_5_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_254;
  reg  conflictPReg_5_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_255;
  reg  conflictPReg_5_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_256;
  reg  conflictPReg_5_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_257;
  reg  conflictPReg_5_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_258;
  reg  conflictPReg_6_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_259;
  reg  conflictPReg_6_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_260;
  reg  conflictPReg_6_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_261;
  reg  conflictPReg_6_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_262;
  reg  conflictPReg_6_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_263;
  reg  conflictPReg_6_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_264;
  reg  conflictPReg_6_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_265;
  reg  conflictPReg_6_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_266;
  reg  conflictPReg_6_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_267;
  reg  conflictPReg_6_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_268;
  reg  conflictPReg_6_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_269;
  reg  conflictPReg_6_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_270;
  reg  conflictPReg_6_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_271;
  reg  conflictPReg_6_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_272;
  reg  conflictPReg_6_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_273;
  reg  conflictPReg_6_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_274;
  reg  conflictPReg_7_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_275;
  reg  conflictPReg_7_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_276;
  reg  conflictPReg_7_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_277;
  reg  conflictPReg_7_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_278;
  reg  conflictPReg_7_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_279;
  reg  conflictPReg_7_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_280;
  reg  conflictPReg_7_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_281;
  reg  conflictPReg_7_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_282;
  reg  conflictPReg_7_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_283;
  reg  conflictPReg_7_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_284;
  reg  conflictPReg_7_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_285;
  reg  conflictPReg_7_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_286;
  reg  conflictPReg_7_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_287;
  reg  conflictPReg_7_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_288;
  reg  conflictPReg_7_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_289;
  reg  conflictPReg_7_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_290;
  reg  conflictPReg_8_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_291;
  reg  conflictPReg_8_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_292;
  reg  conflictPReg_8_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_293;
  reg  conflictPReg_8_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_294;
  reg  conflictPReg_8_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_295;
  reg  conflictPReg_8_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_296;
  reg  conflictPReg_8_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_297;
  reg  conflictPReg_8_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_298;
  reg  conflictPReg_8_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_299;
  reg  conflictPReg_8_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_300;
  reg  conflictPReg_8_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_301;
  reg  conflictPReg_8_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_302;
  reg  conflictPReg_8_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_303;
  reg  conflictPReg_8_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_304;
  reg  conflictPReg_8_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_305;
  reg  conflictPReg_8_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_306;
  reg  conflictPReg_9_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_307;
  reg  conflictPReg_9_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_308;
  reg  conflictPReg_9_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_309;
  reg  conflictPReg_9_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_310;
  reg  conflictPReg_9_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_311;
  reg  conflictPReg_9_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_312;
  reg  conflictPReg_9_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_313;
  reg  conflictPReg_9_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_314;
  reg  conflictPReg_9_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_315;
  reg  conflictPReg_9_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_316;
  reg  conflictPReg_9_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_317;
  reg  conflictPReg_9_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_318;
  reg  conflictPReg_9_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_319;
  reg  conflictPReg_9_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_320;
  reg  conflictPReg_9_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_321;
  reg  conflictPReg_9_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_322;
  reg  conflictPReg_10_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_323;
  reg  conflictPReg_10_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_324;
  reg  conflictPReg_10_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_325;
  reg  conflictPReg_10_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_326;
  reg  conflictPReg_10_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_327;
  reg  conflictPReg_10_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_328;
  reg  conflictPReg_10_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_329;
  reg  conflictPReg_10_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_330;
  reg  conflictPReg_10_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_331;
  reg  conflictPReg_10_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_332;
  reg  conflictPReg_10_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_333;
  reg  conflictPReg_10_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_334;
  reg  conflictPReg_10_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_335;
  reg  conflictPReg_10_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_336;
  reg  conflictPReg_10_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_337;
  reg  conflictPReg_10_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_338;
  reg  conflictPReg_11_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_339;
  reg  conflictPReg_11_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_340;
  reg  conflictPReg_11_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_341;
  reg  conflictPReg_11_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_342;
  reg  conflictPReg_11_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_343;
  reg  conflictPReg_11_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_344;
  reg  conflictPReg_11_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_345;
  reg  conflictPReg_11_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_346;
  reg  conflictPReg_11_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_347;
  reg  conflictPReg_11_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_348;
  reg  conflictPReg_11_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_349;
  reg  conflictPReg_11_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_350;
  reg  conflictPReg_11_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_351;
  reg  conflictPReg_11_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_352;
  reg  conflictPReg_11_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_353;
  reg  conflictPReg_11_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_354;
  reg  conflictPReg_12_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_355;
  reg  conflictPReg_12_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_356;
  reg  conflictPReg_12_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_357;
  reg  conflictPReg_12_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_358;
  reg  conflictPReg_12_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_359;
  reg  conflictPReg_12_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_360;
  reg  conflictPReg_12_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_361;
  reg  conflictPReg_12_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_362;
  reg  conflictPReg_12_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_363;
  reg  conflictPReg_12_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_364;
  reg  conflictPReg_12_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_365;
  reg  conflictPReg_12_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_366;
  reg  conflictPReg_12_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_367;
  reg  conflictPReg_12_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_368;
  reg  conflictPReg_12_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_369;
  reg  conflictPReg_12_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_370;
  reg  conflictPReg_13_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_371;
  reg  conflictPReg_13_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_372;
  reg  conflictPReg_13_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_373;
  reg  conflictPReg_13_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_374;
  reg  conflictPReg_13_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_375;
  reg  conflictPReg_13_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_376;
  reg  conflictPReg_13_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_377;
  reg  conflictPReg_13_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_378;
  reg  conflictPReg_13_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_379;
  reg  conflictPReg_13_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_380;
  reg  conflictPReg_13_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_381;
  reg  conflictPReg_13_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_382;
  reg  conflictPReg_13_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_383;
  reg  conflictPReg_13_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_384;
  reg  conflictPReg_13_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_385;
  reg  conflictPReg_13_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_386;
  reg  conflictPReg_14_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_387;
  reg  conflictPReg_14_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_388;
  reg  conflictPReg_14_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_389;
  reg  conflictPReg_14_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_390;
  reg  conflictPReg_14_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_391;
  reg  conflictPReg_14_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_392;
  reg  conflictPReg_14_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_393;
  reg  conflictPReg_14_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_394;
  reg  conflictPReg_14_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_395;
  reg  conflictPReg_14_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_396;
  reg  conflictPReg_14_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_397;
  reg  conflictPReg_14_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_398;
  reg  conflictPReg_14_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_399;
  reg  conflictPReg_14_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_400;
  reg  conflictPReg_14_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_401;
  reg  conflictPReg_14_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_402;
  reg  conflictPReg_15_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_403;
  reg  conflictPReg_15_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_404;
  reg  conflictPReg_15_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_405;
  reg  conflictPReg_15_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_406;
  reg  conflictPReg_15_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_407;
  reg  conflictPReg_15_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_408;
  reg  conflictPReg_15_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_409;
  reg  conflictPReg_15_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_410;
  reg  conflictPReg_15_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_411;
  reg  conflictPReg_15_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_412;
  reg  conflictPReg_15_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_413;
  reg  conflictPReg_15_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_414;
  reg  conflictPReg_15_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_415;
  reg  conflictPReg_15_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_416;
  reg  conflictPReg_15_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_417;
  reg  conflictPReg_15_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_418;
  wire [7:0] _T_52334; // @[Mux.scala 19:72:@24996.4]
  wire [7:0] _T_52341; // @[Mux.scala 19:72:@25003.4]
  wire [15:0] _T_52342; // @[Mux.scala 19:72:@25004.4]
  wire [15:0] _T_52344; // @[Mux.scala 19:72:@25005.4]
  wire [7:0] _T_52351; // @[Mux.scala 19:72:@25012.4]
  wire [7:0] _T_52358; // @[Mux.scala 19:72:@25019.4]
  wire [15:0] _T_52359; // @[Mux.scala 19:72:@25020.4]
  wire [15:0] _T_52361; // @[Mux.scala 19:72:@25021.4]
  wire [7:0] _T_52368; // @[Mux.scala 19:72:@25028.4]
  wire [7:0] _T_52375; // @[Mux.scala 19:72:@25035.4]
  wire [15:0] _T_52376; // @[Mux.scala 19:72:@25036.4]
  wire [15:0] _T_52378; // @[Mux.scala 19:72:@25037.4]
  wire [7:0] _T_52385; // @[Mux.scala 19:72:@25044.4]
  wire [7:0] _T_52392; // @[Mux.scala 19:72:@25051.4]
  wire [15:0] _T_52393; // @[Mux.scala 19:72:@25052.4]
  wire [15:0] _T_52395; // @[Mux.scala 19:72:@25053.4]
  wire [7:0] _T_52402; // @[Mux.scala 19:72:@25060.4]
  wire [7:0] _T_52409; // @[Mux.scala 19:72:@25067.4]
  wire [15:0] _T_52410; // @[Mux.scala 19:72:@25068.4]
  wire [15:0] _T_52412; // @[Mux.scala 19:72:@25069.4]
  wire [7:0] _T_52419; // @[Mux.scala 19:72:@25076.4]
  wire [7:0] _T_52426; // @[Mux.scala 19:72:@25083.4]
  wire [15:0] _T_52427; // @[Mux.scala 19:72:@25084.4]
  wire [15:0] _T_52429; // @[Mux.scala 19:72:@25085.4]
  wire [7:0] _T_52436; // @[Mux.scala 19:72:@25092.4]
  wire [7:0] _T_52443; // @[Mux.scala 19:72:@25099.4]
  wire [15:0] _T_52444; // @[Mux.scala 19:72:@25100.4]
  wire [15:0] _T_52446; // @[Mux.scala 19:72:@25101.4]
  wire [7:0] _T_52453; // @[Mux.scala 19:72:@25108.4]
  wire [7:0] _T_52460; // @[Mux.scala 19:72:@25115.4]
  wire [15:0] _T_52461; // @[Mux.scala 19:72:@25116.4]
  wire [15:0] _T_52463; // @[Mux.scala 19:72:@25117.4]
  wire [15:0] _T_52478; // @[Mux.scala 19:72:@25132.4]
  wire [15:0] _T_52480; // @[Mux.scala 19:72:@25133.4]
  wire [15:0] _T_52495; // @[Mux.scala 19:72:@25148.4]
  wire [15:0] _T_52497; // @[Mux.scala 19:72:@25149.4]
  wire [15:0] _T_52512; // @[Mux.scala 19:72:@25164.4]
  wire [15:0] _T_52514; // @[Mux.scala 19:72:@25165.4]
  wire [15:0] _T_52529; // @[Mux.scala 19:72:@25180.4]
  wire [15:0] _T_52531; // @[Mux.scala 19:72:@25181.4]
  wire [15:0] _T_52546; // @[Mux.scala 19:72:@25196.4]
  wire [15:0] _T_52548; // @[Mux.scala 19:72:@25197.4]
  wire [15:0] _T_52563; // @[Mux.scala 19:72:@25212.4]
  wire [15:0] _T_52565; // @[Mux.scala 19:72:@25213.4]
  wire [15:0] _T_52580; // @[Mux.scala 19:72:@25228.4]
  wire [15:0] _T_52582; // @[Mux.scala 19:72:@25229.4]
  wire [15:0] _T_52597; // @[Mux.scala 19:72:@25244.4]
  wire [15:0] _T_52599; // @[Mux.scala 19:72:@25245.4]
  wire [15:0] _T_52600; // @[Mux.scala 19:72:@25246.4]
  wire [15:0] _T_52601; // @[Mux.scala 19:72:@25247.4]
  wire [15:0] _T_52602; // @[Mux.scala 19:72:@25248.4]
  wire [15:0] _T_52603; // @[Mux.scala 19:72:@25249.4]
  wire [15:0] _T_52604; // @[Mux.scala 19:72:@25250.4]
  wire [15:0] _T_52605; // @[Mux.scala 19:72:@25251.4]
  wire [15:0] _T_52606; // @[Mux.scala 19:72:@25252.4]
  wire [15:0] _T_52607; // @[Mux.scala 19:72:@25253.4]
  wire [15:0] _T_52608; // @[Mux.scala 19:72:@25254.4]
  wire [15:0] _T_52609; // @[Mux.scala 19:72:@25255.4]
  wire [15:0] _T_52610; // @[Mux.scala 19:72:@25256.4]
  wire [15:0] _T_52611; // @[Mux.scala 19:72:@25257.4]
  wire [15:0] _T_52612; // @[Mux.scala 19:72:@25258.4]
  wire [15:0] _T_52613; // @[Mux.scala 19:72:@25259.4]
  wire [15:0] _T_52614; // @[Mux.scala 19:72:@25260.4]
  wire [7:0] _T_53192; // @[Mux.scala 19:72:@25610.4]
  wire [7:0] _T_53199; // @[Mux.scala 19:72:@25617.4]
  wire [15:0] _T_53200; // @[Mux.scala 19:72:@25618.4]
  wire [15:0] _T_53202; // @[Mux.scala 19:72:@25619.4]
  wire [7:0] _T_53209; // @[Mux.scala 19:72:@25626.4]
  wire [7:0] _T_53216; // @[Mux.scala 19:72:@25633.4]
  wire [15:0] _T_53217; // @[Mux.scala 19:72:@25634.4]
  wire [15:0] _T_53219; // @[Mux.scala 19:72:@25635.4]
  wire [7:0] _T_53226; // @[Mux.scala 19:72:@25642.4]
  wire [7:0] _T_53233; // @[Mux.scala 19:72:@25649.4]
  wire [15:0] _T_53234; // @[Mux.scala 19:72:@25650.4]
  wire [15:0] _T_53236; // @[Mux.scala 19:72:@25651.4]
  wire [7:0] _T_53243; // @[Mux.scala 19:72:@25658.4]
  wire [7:0] _T_53250; // @[Mux.scala 19:72:@25665.4]
  wire [15:0] _T_53251; // @[Mux.scala 19:72:@25666.4]
  wire [15:0] _T_53253; // @[Mux.scala 19:72:@25667.4]
  wire [7:0] _T_53260; // @[Mux.scala 19:72:@25674.4]
  wire [7:0] _T_53267; // @[Mux.scala 19:72:@25681.4]
  wire [15:0] _T_53268; // @[Mux.scala 19:72:@25682.4]
  wire [15:0] _T_53270; // @[Mux.scala 19:72:@25683.4]
  wire [7:0] _T_53277; // @[Mux.scala 19:72:@25690.4]
  wire [7:0] _T_53284; // @[Mux.scala 19:72:@25697.4]
  wire [15:0] _T_53285; // @[Mux.scala 19:72:@25698.4]
  wire [15:0] _T_53287; // @[Mux.scala 19:72:@25699.4]
  wire [7:0] _T_53294; // @[Mux.scala 19:72:@25706.4]
  wire [7:0] _T_53301; // @[Mux.scala 19:72:@25713.4]
  wire [15:0] _T_53302; // @[Mux.scala 19:72:@25714.4]
  wire [15:0] _T_53304; // @[Mux.scala 19:72:@25715.4]
  wire [7:0] _T_53311; // @[Mux.scala 19:72:@25722.4]
  wire [7:0] _T_53318; // @[Mux.scala 19:72:@25729.4]
  wire [15:0] _T_53319; // @[Mux.scala 19:72:@25730.4]
  wire [15:0] _T_53321; // @[Mux.scala 19:72:@25731.4]
  wire [15:0] _T_53336; // @[Mux.scala 19:72:@25746.4]
  wire [15:0] _T_53338; // @[Mux.scala 19:72:@25747.4]
  wire [15:0] _T_53353; // @[Mux.scala 19:72:@25762.4]
  wire [15:0] _T_53355; // @[Mux.scala 19:72:@25763.4]
  wire [15:0] _T_53370; // @[Mux.scala 19:72:@25778.4]
  wire [15:0] _T_53372; // @[Mux.scala 19:72:@25779.4]
  wire [15:0] _T_53387; // @[Mux.scala 19:72:@25794.4]
  wire [15:0] _T_53389; // @[Mux.scala 19:72:@25795.4]
  wire [15:0] _T_53404; // @[Mux.scala 19:72:@25810.4]
  wire [15:0] _T_53406; // @[Mux.scala 19:72:@25811.4]
  wire [15:0] _T_53421; // @[Mux.scala 19:72:@25826.4]
  wire [15:0] _T_53423; // @[Mux.scala 19:72:@25827.4]
  wire [15:0] _T_53438; // @[Mux.scala 19:72:@25842.4]
  wire [15:0] _T_53440; // @[Mux.scala 19:72:@25843.4]
  wire [15:0] _T_53455; // @[Mux.scala 19:72:@25858.4]
  wire [15:0] _T_53457; // @[Mux.scala 19:72:@25859.4]
  wire [15:0] _T_53458; // @[Mux.scala 19:72:@25860.4]
  wire [15:0] _T_53459; // @[Mux.scala 19:72:@25861.4]
  wire [15:0] _T_53460; // @[Mux.scala 19:72:@25862.4]
  wire [15:0] _T_53461; // @[Mux.scala 19:72:@25863.4]
  wire [15:0] _T_53462; // @[Mux.scala 19:72:@25864.4]
  wire [15:0] _T_53463; // @[Mux.scala 19:72:@25865.4]
  wire [15:0] _T_53464; // @[Mux.scala 19:72:@25866.4]
  wire [15:0] _T_53465; // @[Mux.scala 19:72:@25867.4]
  wire [15:0] _T_53466; // @[Mux.scala 19:72:@25868.4]
  wire [15:0] _T_53467; // @[Mux.scala 19:72:@25869.4]
  wire [15:0] _T_53468; // @[Mux.scala 19:72:@25870.4]
  wire [15:0] _T_53469; // @[Mux.scala 19:72:@25871.4]
  wire [15:0] _T_53470; // @[Mux.scala 19:72:@25872.4]
  wire [15:0] _T_53471; // @[Mux.scala 19:72:@25873.4]
  wire [15:0] _T_53472; // @[Mux.scala 19:72:@25874.4]
  wire [7:0] _T_54050; // @[Mux.scala 19:72:@26224.4]
  wire [7:0] _T_54057; // @[Mux.scala 19:72:@26231.4]
  wire [15:0] _T_54058; // @[Mux.scala 19:72:@26232.4]
  wire [15:0] _T_54060; // @[Mux.scala 19:72:@26233.4]
  wire [7:0] _T_54067; // @[Mux.scala 19:72:@26240.4]
  wire [7:0] _T_54074; // @[Mux.scala 19:72:@26247.4]
  wire [15:0] _T_54075; // @[Mux.scala 19:72:@26248.4]
  wire [15:0] _T_54077; // @[Mux.scala 19:72:@26249.4]
  wire [7:0] _T_54084; // @[Mux.scala 19:72:@26256.4]
  wire [7:0] _T_54091; // @[Mux.scala 19:72:@26263.4]
  wire [15:0] _T_54092; // @[Mux.scala 19:72:@26264.4]
  wire [15:0] _T_54094; // @[Mux.scala 19:72:@26265.4]
  wire [7:0] _T_54101; // @[Mux.scala 19:72:@26272.4]
  wire [7:0] _T_54108; // @[Mux.scala 19:72:@26279.4]
  wire [15:0] _T_54109; // @[Mux.scala 19:72:@26280.4]
  wire [15:0] _T_54111; // @[Mux.scala 19:72:@26281.4]
  wire [7:0] _T_54118; // @[Mux.scala 19:72:@26288.4]
  wire [7:0] _T_54125; // @[Mux.scala 19:72:@26295.4]
  wire [15:0] _T_54126; // @[Mux.scala 19:72:@26296.4]
  wire [15:0] _T_54128; // @[Mux.scala 19:72:@26297.4]
  wire [7:0] _T_54135; // @[Mux.scala 19:72:@26304.4]
  wire [7:0] _T_54142; // @[Mux.scala 19:72:@26311.4]
  wire [15:0] _T_54143; // @[Mux.scala 19:72:@26312.4]
  wire [15:0] _T_54145; // @[Mux.scala 19:72:@26313.4]
  wire [7:0] _T_54152; // @[Mux.scala 19:72:@26320.4]
  wire [7:0] _T_54159; // @[Mux.scala 19:72:@26327.4]
  wire [15:0] _T_54160; // @[Mux.scala 19:72:@26328.4]
  wire [15:0] _T_54162; // @[Mux.scala 19:72:@26329.4]
  wire [7:0] _T_54169; // @[Mux.scala 19:72:@26336.4]
  wire [7:0] _T_54176; // @[Mux.scala 19:72:@26343.4]
  wire [15:0] _T_54177; // @[Mux.scala 19:72:@26344.4]
  wire [15:0] _T_54179; // @[Mux.scala 19:72:@26345.4]
  wire [15:0] _T_54194; // @[Mux.scala 19:72:@26360.4]
  wire [15:0] _T_54196; // @[Mux.scala 19:72:@26361.4]
  wire [15:0] _T_54211; // @[Mux.scala 19:72:@26376.4]
  wire [15:0] _T_54213; // @[Mux.scala 19:72:@26377.4]
  wire [15:0] _T_54228; // @[Mux.scala 19:72:@26392.4]
  wire [15:0] _T_54230; // @[Mux.scala 19:72:@26393.4]
  wire [15:0] _T_54245; // @[Mux.scala 19:72:@26408.4]
  wire [15:0] _T_54247; // @[Mux.scala 19:72:@26409.4]
  wire [15:0] _T_54262; // @[Mux.scala 19:72:@26424.4]
  wire [15:0] _T_54264; // @[Mux.scala 19:72:@26425.4]
  wire [15:0] _T_54279; // @[Mux.scala 19:72:@26440.4]
  wire [15:0] _T_54281; // @[Mux.scala 19:72:@26441.4]
  wire [15:0] _T_54296; // @[Mux.scala 19:72:@26456.4]
  wire [15:0] _T_54298; // @[Mux.scala 19:72:@26457.4]
  wire [15:0] _T_54313; // @[Mux.scala 19:72:@26472.4]
  wire [15:0] _T_54315; // @[Mux.scala 19:72:@26473.4]
  wire [15:0] _T_54316; // @[Mux.scala 19:72:@26474.4]
  wire [15:0] _T_54317; // @[Mux.scala 19:72:@26475.4]
  wire [15:0] _T_54318; // @[Mux.scala 19:72:@26476.4]
  wire [15:0] _T_54319; // @[Mux.scala 19:72:@26477.4]
  wire [15:0] _T_54320; // @[Mux.scala 19:72:@26478.4]
  wire [15:0] _T_54321; // @[Mux.scala 19:72:@26479.4]
  wire [15:0] _T_54322; // @[Mux.scala 19:72:@26480.4]
  wire [15:0] _T_54323; // @[Mux.scala 19:72:@26481.4]
  wire [15:0] _T_54324; // @[Mux.scala 19:72:@26482.4]
  wire [15:0] _T_54325; // @[Mux.scala 19:72:@26483.4]
  wire [15:0] _T_54326; // @[Mux.scala 19:72:@26484.4]
  wire [15:0] _T_54327; // @[Mux.scala 19:72:@26485.4]
  wire [15:0] _T_54328; // @[Mux.scala 19:72:@26486.4]
  wire [15:0] _T_54329; // @[Mux.scala 19:72:@26487.4]
  wire [15:0] _T_54330; // @[Mux.scala 19:72:@26488.4]
  wire [7:0] _T_54908; // @[Mux.scala 19:72:@26838.4]
  wire [7:0] _T_54915; // @[Mux.scala 19:72:@26845.4]
  wire [15:0] _T_54916; // @[Mux.scala 19:72:@26846.4]
  wire [15:0] _T_54918; // @[Mux.scala 19:72:@26847.4]
  wire [7:0] _T_54925; // @[Mux.scala 19:72:@26854.4]
  wire [7:0] _T_54932; // @[Mux.scala 19:72:@26861.4]
  wire [15:0] _T_54933; // @[Mux.scala 19:72:@26862.4]
  wire [15:0] _T_54935; // @[Mux.scala 19:72:@26863.4]
  wire [7:0] _T_54942; // @[Mux.scala 19:72:@26870.4]
  wire [7:0] _T_54949; // @[Mux.scala 19:72:@26877.4]
  wire [15:0] _T_54950; // @[Mux.scala 19:72:@26878.4]
  wire [15:0] _T_54952; // @[Mux.scala 19:72:@26879.4]
  wire [7:0] _T_54959; // @[Mux.scala 19:72:@26886.4]
  wire [7:0] _T_54966; // @[Mux.scala 19:72:@26893.4]
  wire [15:0] _T_54967; // @[Mux.scala 19:72:@26894.4]
  wire [15:0] _T_54969; // @[Mux.scala 19:72:@26895.4]
  wire [7:0] _T_54976; // @[Mux.scala 19:72:@26902.4]
  wire [7:0] _T_54983; // @[Mux.scala 19:72:@26909.4]
  wire [15:0] _T_54984; // @[Mux.scala 19:72:@26910.4]
  wire [15:0] _T_54986; // @[Mux.scala 19:72:@26911.4]
  wire [7:0] _T_54993; // @[Mux.scala 19:72:@26918.4]
  wire [7:0] _T_55000; // @[Mux.scala 19:72:@26925.4]
  wire [15:0] _T_55001; // @[Mux.scala 19:72:@26926.4]
  wire [15:0] _T_55003; // @[Mux.scala 19:72:@26927.4]
  wire [7:0] _T_55010; // @[Mux.scala 19:72:@26934.4]
  wire [7:0] _T_55017; // @[Mux.scala 19:72:@26941.4]
  wire [15:0] _T_55018; // @[Mux.scala 19:72:@26942.4]
  wire [15:0] _T_55020; // @[Mux.scala 19:72:@26943.4]
  wire [7:0] _T_55027; // @[Mux.scala 19:72:@26950.4]
  wire [7:0] _T_55034; // @[Mux.scala 19:72:@26957.4]
  wire [15:0] _T_55035; // @[Mux.scala 19:72:@26958.4]
  wire [15:0] _T_55037; // @[Mux.scala 19:72:@26959.4]
  wire [15:0] _T_55052; // @[Mux.scala 19:72:@26974.4]
  wire [15:0] _T_55054; // @[Mux.scala 19:72:@26975.4]
  wire [15:0] _T_55069; // @[Mux.scala 19:72:@26990.4]
  wire [15:0] _T_55071; // @[Mux.scala 19:72:@26991.4]
  wire [15:0] _T_55086; // @[Mux.scala 19:72:@27006.4]
  wire [15:0] _T_55088; // @[Mux.scala 19:72:@27007.4]
  wire [15:0] _T_55103; // @[Mux.scala 19:72:@27022.4]
  wire [15:0] _T_55105; // @[Mux.scala 19:72:@27023.4]
  wire [15:0] _T_55120; // @[Mux.scala 19:72:@27038.4]
  wire [15:0] _T_55122; // @[Mux.scala 19:72:@27039.4]
  wire [15:0] _T_55137; // @[Mux.scala 19:72:@27054.4]
  wire [15:0] _T_55139; // @[Mux.scala 19:72:@27055.4]
  wire [15:0] _T_55154; // @[Mux.scala 19:72:@27070.4]
  wire [15:0] _T_55156; // @[Mux.scala 19:72:@27071.4]
  wire [15:0] _T_55171; // @[Mux.scala 19:72:@27086.4]
  wire [15:0] _T_55173; // @[Mux.scala 19:72:@27087.4]
  wire [15:0] _T_55174; // @[Mux.scala 19:72:@27088.4]
  wire [15:0] _T_55175; // @[Mux.scala 19:72:@27089.4]
  wire [15:0] _T_55176; // @[Mux.scala 19:72:@27090.4]
  wire [15:0] _T_55177; // @[Mux.scala 19:72:@27091.4]
  wire [15:0] _T_55178; // @[Mux.scala 19:72:@27092.4]
  wire [15:0] _T_55179; // @[Mux.scala 19:72:@27093.4]
  wire [15:0] _T_55180; // @[Mux.scala 19:72:@27094.4]
  wire [15:0] _T_55181; // @[Mux.scala 19:72:@27095.4]
  wire [15:0] _T_55182; // @[Mux.scala 19:72:@27096.4]
  wire [15:0] _T_55183; // @[Mux.scala 19:72:@27097.4]
  wire [15:0] _T_55184; // @[Mux.scala 19:72:@27098.4]
  wire [15:0] _T_55185; // @[Mux.scala 19:72:@27099.4]
  wire [15:0] _T_55186; // @[Mux.scala 19:72:@27100.4]
  wire [15:0] _T_55187; // @[Mux.scala 19:72:@27101.4]
  wire [15:0] _T_55188; // @[Mux.scala 19:72:@27102.4]
  wire [7:0] _T_55766; // @[Mux.scala 19:72:@27452.4]
  wire [7:0] _T_55773; // @[Mux.scala 19:72:@27459.4]
  wire [15:0] _T_55774; // @[Mux.scala 19:72:@27460.4]
  wire [15:0] _T_55776; // @[Mux.scala 19:72:@27461.4]
  wire [7:0] _T_55783; // @[Mux.scala 19:72:@27468.4]
  wire [7:0] _T_55790; // @[Mux.scala 19:72:@27475.4]
  wire [15:0] _T_55791; // @[Mux.scala 19:72:@27476.4]
  wire [15:0] _T_55793; // @[Mux.scala 19:72:@27477.4]
  wire [7:0] _T_55800; // @[Mux.scala 19:72:@27484.4]
  wire [7:0] _T_55807; // @[Mux.scala 19:72:@27491.4]
  wire [15:0] _T_55808; // @[Mux.scala 19:72:@27492.4]
  wire [15:0] _T_55810; // @[Mux.scala 19:72:@27493.4]
  wire [7:0] _T_55817; // @[Mux.scala 19:72:@27500.4]
  wire [7:0] _T_55824; // @[Mux.scala 19:72:@27507.4]
  wire [15:0] _T_55825; // @[Mux.scala 19:72:@27508.4]
  wire [15:0] _T_55827; // @[Mux.scala 19:72:@27509.4]
  wire [7:0] _T_55834; // @[Mux.scala 19:72:@27516.4]
  wire [7:0] _T_55841; // @[Mux.scala 19:72:@27523.4]
  wire [15:0] _T_55842; // @[Mux.scala 19:72:@27524.4]
  wire [15:0] _T_55844; // @[Mux.scala 19:72:@27525.4]
  wire [7:0] _T_55851; // @[Mux.scala 19:72:@27532.4]
  wire [7:0] _T_55858; // @[Mux.scala 19:72:@27539.4]
  wire [15:0] _T_55859; // @[Mux.scala 19:72:@27540.4]
  wire [15:0] _T_55861; // @[Mux.scala 19:72:@27541.4]
  wire [7:0] _T_55868; // @[Mux.scala 19:72:@27548.4]
  wire [7:0] _T_55875; // @[Mux.scala 19:72:@27555.4]
  wire [15:0] _T_55876; // @[Mux.scala 19:72:@27556.4]
  wire [15:0] _T_55878; // @[Mux.scala 19:72:@27557.4]
  wire [7:0] _T_55885; // @[Mux.scala 19:72:@27564.4]
  wire [7:0] _T_55892; // @[Mux.scala 19:72:@27571.4]
  wire [15:0] _T_55893; // @[Mux.scala 19:72:@27572.4]
  wire [15:0] _T_55895; // @[Mux.scala 19:72:@27573.4]
  wire [15:0] _T_55910; // @[Mux.scala 19:72:@27588.4]
  wire [15:0] _T_55912; // @[Mux.scala 19:72:@27589.4]
  wire [15:0] _T_55927; // @[Mux.scala 19:72:@27604.4]
  wire [15:0] _T_55929; // @[Mux.scala 19:72:@27605.4]
  wire [15:0] _T_55944; // @[Mux.scala 19:72:@27620.4]
  wire [15:0] _T_55946; // @[Mux.scala 19:72:@27621.4]
  wire [15:0] _T_55961; // @[Mux.scala 19:72:@27636.4]
  wire [15:0] _T_55963; // @[Mux.scala 19:72:@27637.4]
  wire [15:0] _T_55978; // @[Mux.scala 19:72:@27652.4]
  wire [15:0] _T_55980; // @[Mux.scala 19:72:@27653.4]
  wire [15:0] _T_55995; // @[Mux.scala 19:72:@27668.4]
  wire [15:0] _T_55997; // @[Mux.scala 19:72:@27669.4]
  wire [15:0] _T_56012; // @[Mux.scala 19:72:@27684.4]
  wire [15:0] _T_56014; // @[Mux.scala 19:72:@27685.4]
  wire [15:0] _T_56029; // @[Mux.scala 19:72:@27700.4]
  wire [15:0] _T_56031; // @[Mux.scala 19:72:@27701.4]
  wire [15:0] _T_56032; // @[Mux.scala 19:72:@27702.4]
  wire [15:0] _T_56033; // @[Mux.scala 19:72:@27703.4]
  wire [15:0] _T_56034; // @[Mux.scala 19:72:@27704.4]
  wire [15:0] _T_56035; // @[Mux.scala 19:72:@27705.4]
  wire [15:0] _T_56036; // @[Mux.scala 19:72:@27706.4]
  wire [15:0] _T_56037; // @[Mux.scala 19:72:@27707.4]
  wire [15:0] _T_56038; // @[Mux.scala 19:72:@27708.4]
  wire [15:0] _T_56039; // @[Mux.scala 19:72:@27709.4]
  wire [15:0] _T_56040; // @[Mux.scala 19:72:@27710.4]
  wire [15:0] _T_56041; // @[Mux.scala 19:72:@27711.4]
  wire [15:0] _T_56042; // @[Mux.scala 19:72:@27712.4]
  wire [15:0] _T_56043; // @[Mux.scala 19:72:@27713.4]
  wire [15:0] _T_56044; // @[Mux.scala 19:72:@27714.4]
  wire [15:0] _T_56045; // @[Mux.scala 19:72:@27715.4]
  wire [15:0] _T_56046; // @[Mux.scala 19:72:@27716.4]
  wire [7:0] _T_56624; // @[Mux.scala 19:72:@28066.4]
  wire [7:0] _T_56631; // @[Mux.scala 19:72:@28073.4]
  wire [15:0] _T_56632; // @[Mux.scala 19:72:@28074.4]
  wire [15:0] _T_56634; // @[Mux.scala 19:72:@28075.4]
  wire [7:0] _T_56641; // @[Mux.scala 19:72:@28082.4]
  wire [7:0] _T_56648; // @[Mux.scala 19:72:@28089.4]
  wire [15:0] _T_56649; // @[Mux.scala 19:72:@28090.4]
  wire [15:0] _T_56651; // @[Mux.scala 19:72:@28091.4]
  wire [7:0] _T_56658; // @[Mux.scala 19:72:@28098.4]
  wire [7:0] _T_56665; // @[Mux.scala 19:72:@28105.4]
  wire [15:0] _T_56666; // @[Mux.scala 19:72:@28106.4]
  wire [15:0] _T_56668; // @[Mux.scala 19:72:@28107.4]
  wire [7:0] _T_56675; // @[Mux.scala 19:72:@28114.4]
  wire [7:0] _T_56682; // @[Mux.scala 19:72:@28121.4]
  wire [15:0] _T_56683; // @[Mux.scala 19:72:@28122.4]
  wire [15:0] _T_56685; // @[Mux.scala 19:72:@28123.4]
  wire [7:0] _T_56692; // @[Mux.scala 19:72:@28130.4]
  wire [7:0] _T_56699; // @[Mux.scala 19:72:@28137.4]
  wire [15:0] _T_56700; // @[Mux.scala 19:72:@28138.4]
  wire [15:0] _T_56702; // @[Mux.scala 19:72:@28139.4]
  wire [7:0] _T_56709; // @[Mux.scala 19:72:@28146.4]
  wire [7:0] _T_56716; // @[Mux.scala 19:72:@28153.4]
  wire [15:0] _T_56717; // @[Mux.scala 19:72:@28154.4]
  wire [15:0] _T_56719; // @[Mux.scala 19:72:@28155.4]
  wire [7:0] _T_56726; // @[Mux.scala 19:72:@28162.4]
  wire [7:0] _T_56733; // @[Mux.scala 19:72:@28169.4]
  wire [15:0] _T_56734; // @[Mux.scala 19:72:@28170.4]
  wire [15:0] _T_56736; // @[Mux.scala 19:72:@28171.4]
  wire [7:0] _T_56743; // @[Mux.scala 19:72:@28178.4]
  wire [7:0] _T_56750; // @[Mux.scala 19:72:@28185.4]
  wire [15:0] _T_56751; // @[Mux.scala 19:72:@28186.4]
  wire [15:0] _T_56753; // @[Mux.scala 19:72:@28187.4]
  wire [15:0] _T_56768; // @[Mux.scala 19:72:@28202.4]
  wire [15:0] _T_56770; // @[Mux.scala 19:72:@28203.4]
  wire [15:0] _T_56785; // @[Mux.scala 19:72:@28218.4]
  wire [15:0] _T_56787; // @[Mux.scala 19:72:@28219.4]
  wire [15:0] _T_56802; // @[Mux.scala 19:72:@28234.4]
  wire [15:0] _T_56804; // @[Mux.scala 19:72:@28235.4]
  wire [15:0] _T_56819; // @[Mux.scala 19:72:@28250.4]
  wire [15:0] _T_56821; // @[Mux.scala 19:72:@28251.4]
  wire [15:0] _T_56836; // @[Mux.scala 19:72:@28266.4]
  wire [15:0] _T_56838; // @[Mux.scala 19:72:@28267.4]
  wire [15:0] _T_56853; // @[Mux.scala 19:72:@28282.4]
  wire [15:0] _T_56855; // @[Mux.scala 19:72:@28283.4]
  wire [15:0] _T_56870; // @[Mux.scala 19:72:@28298.4]
  wire [15:0] _T_56872; // @[Mux.scala 19:72:@28299.4]
  wire [15:0] _T_56887; // @[Mux.scala 19:72:@28314.4]
  wire [15:0] _T_56889; // @[Mux.scala 19:72:@28315.4]
  wire [15:0] _T_56890; // @[Mux.scala 19:72:@28316.4]
  wire [15:0] _T_56891; // @[Mux.scala 19:72:@28317.4]
  wire [15:0] _T_56892; // @[Mux.scala 19:72:@28318.4]
  wire [15:0] _T_56893; // @[Mux.scala 19:72:@28319.4]
  wire [15:0] _T_56894; // @[Mux.scala 19:72:@28320.4]
  wire [15:0] _T_56895; // @[Mux.scala 19:72:@28321.4]
  wire [15:0] _T_56896; // @[Mux.scala 19:72:@28322.4]
  wire [15:0] _T_56897; // @[Mux.scala 19:72:@28323.4]
  wire [15:0] _T_56898; // @[Mux.scala 19:72:@28324.4]
  wire [15:0] _T_56899; // @[Mux.scala 19:72:@28325.4]
  wire [15:0] _T_56900; // @[Mux.scala 19:72:@28326.4]
  wire [15:0] _T_56901; // @[Mux.scala 19:72:@28327.4]
  wire [15:0] _T_56902; // @[Mux.scala 19:72:@28328.4]
  wire [15:0] _T_56903; // @[Mux.scala 19:72:@28329.4]
  wire [15:0] _T_56904; // @[Mux.scala 19:72:@28330.4]
  wire [7:0] _T_57482; // @[Mux.scala 19:72:@28680.4]
  wire [7:0] _T_57489; // @[Mux.scala 19:72:@28687.4]
  wire [15:0] _T_57490; // @[Mux.scala 19:72:@28688.4]
  wire [15:0] _T_57492; // @[Mux.scala 19:72:@28689.4]
  wire [7:0] _T_57499; // @[Mux.scala 19:72:@28696.4]
  wire [7:0] _T_57506; // @[Mux.scala 19:72:@28703.4]
  wire [15:0] _T_57507; // @[Mux.scala 19:72:@28704.4]
  wire [15:0] _T_57509; // @[Mux.scala 19:72:@28705.4]
  wire [7:0] _T_57516; // @[Mux.scala 19:72:@28712.4]
  wire [7:0] _T_57523; // @[Mux.scala 19:72:@28719.4]
  wire [15:0] _T_57524; // @[Mux.scala 19:72:@28720.4]
  wire [15:0] _T_57526; // @[Mux.scala 19:72:@28721.4]
  wire [7:0] _T_57533; // @[Mux.scala 19:72:@28728.4]
  wire [7:0] _T_57540; // @[Mux.scala 19:72:@28735.4]
  wire [15:0] _T_57541; // @[Mux.scala 19:72:@28736.4]
  wire [15:0] _T_57543; // @[Mux.scala 19:72:@28737.4]
  wire [7:0] _T_57550; // @[Mux.scala 19:72:@28744.4]
  wire [7:0] _T_57557; // @[Mux.scala 19:72:@28751.4]
  wire [15:0] _T_57558; // @[Mux.scala 19:72:@28752.4]
  wire [15:0] _T_57560; // @[Mux.scala 19:72:@28753.4]
  wire [7:0] _T_57567; // @[Mux.scala 19:72:@28760.4]
  wire [7:0] _T_57574; // @[Mux.scala 19:72:@28767.4]
  wire [15:0] _T_57575; // @[Mux.scala 19:72:@28768.4]
  wire [15:0] _T_57577; // @[Mux.scala 19:72:@28769.4]
  wire [7:0] _T_57584; // @[Mux.scala 19:72:@28776.4]
  wire [7:0] _T_57591; // @[Mux.scala 19:72:@28783.4]
  wire [15:0] _T_57592; // @[Mux.scala 19:72:@28784.4]
  wire [15:0] _T_57594; // @[Mux.scala 19:72:@28785.4]
  wire [7:0] _T_57601; // @[Mux.scala 19:72:@28792.4]
  wire [7:0] _T_57608; // @[Mux.scala 19:72:@28799.4]
  wire [15:0] _T_57609; // @[Mux.scala 19:72:@28800.4]
  wire [15:0] _T_57611; // @[Mux.scala 19:72:@28801.4]
  wire [15:0] _T_57626; // @[Mux.scala 19:72:@28816.4]
  wire [15:0] _T_57628; // @[Mux.scala 19:72:@28817.4]
  wire [15:0] _T_57643; // @[Mux.scala 19:72:@28832.4]
  wire [15:0] _T_57645; // @[Mux.scala 19:72:@28833.4]
  wire [15:0] _T_57660; // @[Mux.scala 19:72:@28848.4]
  wire [15:0] _T_57662; // @[Mux.scala 19:72:@28849.4]
  wire [15:0] _T_57677; // @[Mux.scala 19:72:@28864.4]
  wire [15:0] _T_57679; // @[Mux.scala 19:72:@28865.4]
  wire [15:0] _T_57694; // @[Mux.scala 19:72:@28880.4]
  wire [15:0] _T_57696; // @[Mux.scala 19:72:@28881.4]
  wire [15:0] _T_57711; // @[Mux.scala 19:72:@28896.4]
  wire [15:0] _T_57713; // @[Mux.scala 19:72:@28897.4]
  wire [15:0] _T_57728; // @[Mux.scala 19:72:@28912.4]
  wire [15:0] _T_57730; // @[Mux.scala 19:72:@28913.4]
  wire [15:0] _T_57745; // @[Mux.scala 19:72:@28928.4]
  wire [15:0] _T_57747; // @[Mux.scala 19:72:@28929.4]
  wire [15:0] _T_57748; // @[Mux.scala 19:72:@28930.4]
  wire [15:0] _T_57749; // @[Mux.scala 19:72:@28931.4]
  wire [15:0] _T_57750; // @[Mux.scala 19:72:@28932.4]
  wire [15:0] _T_57751; // @[Mux.scala 19:72:@28933.4]
  wire [15:0] _T_57752; // @[Mux.scala 19:72:@28934.4]
  wire [15:0] _T_57753; // @[Mux.scala 19:72:@28935.4]
  wire [15:0] _T_57754; // @[Mux.scala 19:72:@28936.4]
  wire [15:0] _T_57755; // @[Mux.scala 19:72:@28937.4]
  wire [15:0] _T_57756; // @[Mux.scala 19:72:@28938.4]
  wire [15:0] _T_57757; // @[Mux.scala 19:72:@28939.4]
  wire [15:0] _T_57758; // @[Mux.scala 19:72:@28940.4]
  wire [15:0] _T_57759; // @[Mux.scala 19:72:@28941.4]
  wire [15:0] _T_57760; // @[Mux.scala 19:72:@28942.4]
  wire [15:0] _T_57761; // @[Mux.scala 19:72:@28943.4]
  wire [15:0] _T_57762; // @[Mux.scala 19:72:@28944.4]
  wire [7:0] _T_58340; // @[Mux.scala 19:72:@29294.4]
  wire [7:0] _T_58347; // @[Mux.scala 19:72:@29301.4]
  wire [15:0] _T_58348; // @[Mux.scala 19:72:@29302.4]
  wire [15:0] _T_58350; // @[Mux.scala 19:72:@29303.4]
  wire [7:0] _T_58357; // @[Mux.scala 19:72:@29310.4]
  wire [7:0] _T_58364; // @[Mux.scala 19:72:@29317.4]
  wire [15:0] _T_58365; // @[Mux.scala 19:72:@29318.4]
  wire [15:0] _T_58367; // @[Mux.scala 19:72:@29319.4]
  wire [7:0] _T_58374; // @[Mux.scala 19:72:@29326.4]
  wire [7:0] _T_58381; // @[Mux.scala 19:72:@29333.4]
  wire [15:0] _T_58382; // @[Mux.scala 19:72:@29334.4]
  wire [15:0] _T_58384; // @[Mux.scala 19:72:@29335.4]
  wire [7:0] _T_58391; // @[Mux.scala 19:72:@29342.4]
  wire [7:0] _T_58398; // @[Mux.scala 19:72:@29349.4]
  wire [15:0] _T_58399; // @[Mux.scala 19:72:@29350.4]
  wire [15:0] _T_58401; // @[Mux.scala 19:72:@29351.4]
  wire [7:0] _T_58408; // @[Mux.scala 19:72:@29358.4]
  wire [7:0] _T_58415; // @[Mux.scala 19:72:@29365.4]
  wire [15:0] _T_58416; // @[Mux.scala 19:72:@29366.4]
  wire [15:0] _T_58418; // @[Mux.scala 19:72:@29367.4]
  wire [7:0] _T_58425; // @[Mux.scala 19:72:@29374.4]
  wire [7:0] _T_58432; // @[Mux.scala 19:72:@29381.4]
  wire [15:0] _T_58433; // @[Mux.scala 19:72:@29382.4]
  wire [15:0] _T_58435; // @[Mux.scala 19:72:@29383.4]
  wire [7:0] _T_58442; // @[Mux.scala 19:72:@29390.4]
  wire [7:0] _T_58449; // @[Mux.scala 19:72:@29397.4]
  wire [15:0] _T_58450; // @[Mux.scala 19:72:@29398.4]
  wire [15:0] _T_58452; // @[Mux.scala 19:72:@29399.4]
  wire [7:0] _T_58459; // @[Mux.scala 19:72:@29406.4]
  wire [7:0] _T_58466; // @[Mux.scala 19:72:@29413.4]
  wire [15:0] _T_58467; // @[Mux.scala 19:72:@29414.4]
  wire [15:0] _T_58469; // @[Mux.scala 19:72:@29415.4]
  wire [15:0] _T_58484; // @[Mux.scala 19:72:@29430.4]
  wire [15:0] _T_58486; // @[Mux.scala 19:72:@29431.4]
  wire [15:0] _T_58501; // @[Mux.scala 19:72:@29446.4]
  wire [15:0] _T_58503; // @[Mux.scala 19:72:@29447.4]
  wire [15:0] _T_58518; // @[Mux.scala 19:72:@29462.4]
  wire [15:0] _T_58520; // @[Mux.scala 19:72:@29463.4]
  wire [15:0] _T_58535; // @[Mux.scala 19:72:@29478.4]
  wire [15:0] _T_58537; // @[Mux.scala 19:72:@29479.4]
  wire [15:0] _T_58552; // @[Mux.scala 19:72:@29494.4]
  wire [15:0] _T_58554; // @[Mux.scala 19:72:@29495.4]
  wire [15:0] _T_58569; // @[Mux.scala 19:72:@29510.4]
  wire [15:0] _T_58571; // @[Mux.scala 19:72:@29511.4]
  wire [15:0] _T_58586; // @[Mux.scala 19:72:@29526.4]
  wire [15:0] _T_58588; // @[Mux.scala 19:72:@29527.4]
  wire [15:0] _T_58603; // @[Mux.scala 19:72:@29542.4]
  wire [15:0] _T_58605; // @[Mux.scala 19:72:@29543.4]
  wire [15:0] _T_58606; // @[Mux.scala 19:72:@29544.4]
  wire [15:0] _T_58607; // @[Mux.scala 19:72:@29545.4]
  wire [15:0] _T_58608; // @[Mux.scala 19:72:@29546.4]
  wire [15:0] _T_58609; // @[Mux.scala 19:72:@29547.4]
  wire [15:0] _T_58610; // @[Mux.scala 19:72:@29548.4]
  wire [15:0] _T_58611; // @[Mux.scala 19:72:@29549.4]
  wire [15:0] _T_58612; // @[Mux.scala 19:72:@29550.4]
  wire [15:0] _T_58613; // @[Mux.scala 19:72:@29551.4]
  wire [15:0] _T_58614; // @[Mux.scala 19:72:@29552.4]
  wire [15:0] _T_58615; // @[Mux.scala 19:72:@29553.4]
  wire [15:0] _T_58616; // @[Mux.scala 19:72:@29554.4]
  wire [15:0] _T_58617; // @[Mux.scala 19:72:@29555.4]
  wire [15:0] _T_58618; // @[Mux.scala 19:72:@29556.4]
  wire [15:0] _T_58619; // @[Mux.scala 19:72:@29557.4]
  wire [15:0] _T_58620; // @[Mux.scala 19:72:@29558.4]
  wire [7:0] _T_59198; // @[Mux.scala 19:72:@29908.4]
  wire [7:0] _T_59205; // @[Mux.scala 19:72:@29915.4]
  wire [15:0] _T_59206; // @[Mux.scala 19:72:@29916.4]
  wire [15:0] _T_59208; // @[Mux.scala 19:72:@29917.4]
  wire [7:0] _T_59215; // @[Mux.scala 19:72:@29924.4]
  wire [7:0] _T_59222; // @[Mux.scala 19:72:@29931.4]
  wire [15:0] _T_59223; // @[Mux.scala 19:72:@29932.4]
  wire [15:0] _T_59225; // @[Mux.scala 19:72:@29933.4]
  wire [7:0] _T_59232; // @[Mux.scala 19:72:@29940.4]
  wire [7:0] _T_59239; // @[Mux.scala 19:72:@29947.4]
  wire [15:0] _T_59240; // @[Mux.scala 19:72:@29948.4]
  wire [15:0] _T_59242; // @[Mux.scala 19:72:@29949.4]
  wire [7:0] _T_59249; // @[Mux.scala 19:72:@29956.4]
  wire [7:0] _T_59256; // @[Mux.scala 19:72:@29963.4]
  wire [15:0] _T_59257; // @[Mux.scala 19:72:@29964.4]
  wire [15:0] _T_59259; // @[Mux.scala 19:72:@29965.4]
  wire [7:0] _T_59266; // @[Mux.scala 19:72:@29972.4]
  wire [7:0] _T_59273; // @[Mux.scala 19:72:@29979.4]
  wire [15:0] _T_59274; // @[Mux.scala 19:72:@29980.4]
  wire [15:0] _T_59276; // @[Mux.scala 19:72:@29981.4]
  wire [7:0] _T_59283; // @[Mux.scala 19:72:@29988.4]
  wire [7:0] _T_59290; // @[Mux.scala 19:72:@29995.4]
  wire [15:0] _T_59291; // @[Mux.scala 19:72:@29996.4]
  wire [15:0] _T_59293; // @[Mux.scala 19:72:@29997.4]
  wire [7:0] _T_59300; // @[Mux.scala 19:72:@30004.4]
  wire [7:0] _T_59307; // @[Mux.scala 19:72:@30011.4]
  wire [15:0] _T_59308; // @[Mux.scala 19:72:@30012.4]
  wire [15:0] _T_59310; // @[Mux.scala 19:72:@30013.4]
  wire [7:0] _T_59317; // @[Mux.scala 19:72:@30020.4]
  wire [7:0] _T_59324; // @[Mux.scala 19:72:@30027.4]
  wire [15:0] _T_59325; // @[Mux.scala 19:72:@30028.4]
  wire [15:0] _T_59327; // @[Mux.scala 19:72:@30029.4]
  wire [15:0] _T_59342; // @[Mux.scala 19:72:@30044.4]
  wire [15:0] _T_59344; // @[Mux.scala 19:72:@30045.4]
  wire [15:0] _T_59359; // @[Mux.scala 19:72:@30060.4]
  wire [15:0] _T_59361; // @[Mux.scala 19:72:@30061.4]
  wire [15:0] _T_59376; // @[Mux.scala 19:72:@30076.4]
  wire [15:0] _T_59378; // @[Mux.scala 19:72:@30077.4]
  wire [15:0] _T_59393; // @[Mux.scala 19:72:@30092.4]
  wire [15:0] _T_59395; // @[Mux.scala 19:72:@30093.4]
  wire [15:0] _T_59410; // @[Mux.scala 19:72:@30108.4]
  wire [15:0] _T_59412; // @[Mux.scala 19:72:@30109.4]
  wire [15:0] _T_59427; // @[Mux.scala 19:72:@30124.4]
  wire [15:0] _T_59429; // @[Mux.scala 19:72:@30125.4]
  wire [15:0] _T_59444; // @[Mux.scala 19:72:@30140.4]
  wire [15:0] _T_59446; // @[Mux.scala 19:72:@30141.4]
  wire [15:0] _T_59461; // @[Mux.scala 19:72:@30156.4]
  wire [15:0] _T_59463; // @[Mux.scala 19:72:@30157.4]
  wire [15:0] _T_59464; // @[Mux.scala 19:72:@30158.4]
  wire [15:0] _T_59465; // @[Mux.scala 19:72:@30159.4]
  wire [15:0] _T_59466; // @[Mux.scala 19:72:@30160.4]
  wire [15:0] _T_59467; // @[Mux.scala 19:72:@30161.4]
  wire [15:0] _T_59468; // @[Mux.scala 19:72:@30162.4]
  wire [15:0] _T_59469; // @[Mux.scala 19:72:@30163.4]
  wire [15:0] _T_59470; // @[Mux.scala 19:72:@30164.4]
  wire [15:0] _T_59471; // @[Mux.scala 19:72:@30165.4]
  wire [15:0] _T_59472; // @[Mux.scala 19:72:@30166.4]
  wire [15:0] _T_59473; // @[Mux.scala 19:72:@30167.4]
  wire [15:0] _T_59474; // @[Mux.scala 19:72:@30168.4]
  wire [15:0] _T_59475; // @[Mux.scala 19:72:@30169.4]
  wire [15:0] _T_59476; // @[Mux.scala 19:72:@30170.4]
  wire [15:0] _T_59477; // @[Mux.scala 19:72:@30171.4]
  wire [15:0] _T_59478; // @[Mux.scala 19:72:@30172.4]
  wire [7:0] _T_60056; // @[Mux.scala 19:72:@30522.4]
  wire [7:0] _T_60063; // @[Mux.scala 19:72:@30529.4]
  wire [15:0] _T_60064; // @[Mux.scala 19:72:@30530.4]
  wire [15:0] _T_60066; // @[Mux.scala 19:72:@30531.4]
  wire [7:0] _T_60073; // @[Mux.scala 19:72:@30538.4]
  wire [7:0] _T_60080; // @[Mux.scala 19:72:@30545.4]
  wire [15:0] _T_60081; // @[Mux.scala 19:72:@30546.4]
  wire [15:0] _T_60083; // @[Mux.scala 19:72:@30547.4]
  wire [7:0] _T_60090; // @[Mux.scala 19:72:@30554.4]
  wire [7:0] _T_60097; // @[Mux.scala 19:72:@30561.4]
  wire [15:0] _T_60098; // @[Mux.scala 19:72:@30562.4]
  wire [15:0] _T_60100; // @[Mux.scala 19:72:@30563.4]
  wire [7:0] _T_60107; // @[Mux.scala 19:72:@30570.4]
  wire [7:0] _T_60114; // @[Mux.scala 19:72:@30577.4]
  wire [15:0] _T_60115; // @[Mux.scala 19:72:@30578.4]
  wire [15:0] _T_60117; // @[Mux.scala 19:72:@30579.4]
  wire [7:0] _T_60124; // @[Mux.scala 19:72:@30586.4]
  wire [7:0] _T_60131; // @[Mux.scala 19:72:@30593.4]
  wire [15:0] _T_60132; // @[Mux.scala 19:72:@30594.4]
  wire [15:0] _T_60134; // @[Mux.scala 19:72:@30595.4]
  wire [7:0] _T_60141; // @[Mux.scala 19:72:@30602.4]
  wire [7:0] _T_60148; // @[Mux.scala 19:72:@30609.4]
  wire [15:0] _T_60149; // @[Mux.scala 19:72:@30610.4]
  wire [15:0] _T_60151; // @[Mux.scala 19:72:@30611.4]
  wire [7:0] _T_60158; // @[Mux.scala 19:72:@30618.4]
  wire [7:0] _T_60165; // @[Mux.scala 19:72:@30625.4]
  wire [15:0] _T_60166; // @[Mux.scala 19:72:@30626.4]
  wire [15:0] _T_60168; // @[Mux.scala 19:72:@30627.4]
  wire [7:0] _T_60175; // @[Mux.scala 19:72:@30634.4]
  wire [7:0] _T_60182; // @[Mux.scala 19:72:@30641.4]
  wire [15:0] _T_60183; // @[Mux.scala 19:72:@30642.4]
  wire [15:0] _T_60185; // @[Mux.scala 19:72:@30643.4]
  wire [15:0] _T_60200; // @[Mux.scala 19:72:@30658.4]
  wire [15:0] _T_60202; // @[Mux.scala 19:72:@30659.4]
  wire [15:0] _T_60217; // @[Mux.scala 19:72:@30674.4]
  wire [15:0] _T_60219; // @[Mux.scala 19:72:@30675.4]
  wire [15:0] _T_60234; // @[Mux.scala 19:72:@30690.4]
  wire [15:0] _T_60236; // @[Mux.scala 19:72:@30691.4]
  wire [15:0] _T_60251; // @[Mux.scala 19:72:@30706.4]
  wire [15:0] _T_60253; // @[Mux.scala 19:72:@30707.4]
  wire [15:0] _T_60268; // @[Mux.scala 19:72:@30722.4]
  wire [15:0] _T_60270; // @[Mux.scala 19:72:@30723.4]
  wire [15:0] _T_60285; // @[Mux.scala 19:72:@30738.4]
  wire [15:0] _T_60287; // @[Mux.scala 19:72:@30739.4]
  wire [15:0] _T_60302; // @[Mux.scala 19:72:@30754.4]
  wire [15:0] _T_60304; // @[Mux.scala 19:72:@30755.4]
  wire [15:0] _T_60319; // @[Mux.scala 19:72:@30770.4]
  wire [15:0] _T_60321; // @[Mux.scala 19:72:@30771.4]
  wire [15:0] _T_60322; // @[Mux.scala 19:72:@30772.4]
  wire [15:0] _T_60323; // @[Mux.scala 19:72:@30773.4]
  wire [15:0] _T_60324; // @[Mux.scala 19:72:@30774.4]
  wire [15:0] _T_60325; // @[Mux.scala 19:72:@30775.4]
  wire [15:0] _T_60326; // @[Mux.scala 19:72:@30776.4]
  wire [15:0] _T_60327; // @[Mux.scala 19:72:@30777.4]
  wire [15:0] _T_60328; // @[Mux.scala 19:72:@30778.4]
  wire [15:0] _T_60329; // @[Mux.scala 19:72:@30779.4]
  wire [15:0] _T_60330; // @[Mux.scala 19:72:@30780.4]
  wire [15:0] _T_60331; // @[Mux.scala 19:72:@30781.4]
  wire [15:0] _T_60332; // @[Mux.scala 19:72:@30782.4]
  wire [15:0] _T_60333; // @[Mux.scala 19:72:@30783.4]
  wire [15:0] _T_60334; // @[Mux.scala 19:72:@30784.4]
  wire [15:0] _T_60335; // @[Mux.scala 19:72:@30785.4]
  wire [15:0] _T_60336; // @[Mux.scala 19:72:@30786.4]
  wire [7:0] _T_60914; // @[Mux.scala 19:72:@31136.4]
  wire [7:0] _T_60921; // @[Mux.scala 19:72:@31143.4]
  wire [15:0] _T_60922; // @[Mux.scala 19:72:@31144.4]
  wire [15:0] _T_60924; // @[Mux.scala 19:72:@31145.4]
  wire [7:0] _T_60931; // @[Mux.scala 19:72:@31152.4]
  wire [7:0] _T_60938; // @[Mux.scala 19:72:@31159.4]
  wire [15:0] _T_60939; // @[Mux.scala 19:72:@31160.4]
  wire [15:0] _T_60941; // @[Mux.scala 19:72:@31161.4]
  wire [7:0] _T_60948; // @[Mux.scala 19:72:@31168.4]
  wire [7:0] _T_60955; // @[Mux.scala 19:72:@31175.4]
  wire [15:0] _T_60956; // @[Mux.scala 19:72:@31176.4]
  wire [15:0] _T_60958; // @[Mux.scala 19:72:@31177.4]
  wire [7:0] _T_60965; // @[Mux.scala 19:72:@31184.4]
  wire [7:0] _T_60972; // @[Mux.scala 19:72:@31191.4]
  wire [15:0] _T_60973; // @[Mux.scala 19:72:@31192.4]
  wire [15:0] _T_60975; // @[Mux.scala 19:72:@31193.4]
  wire [7:0] _T_60982; // @[Mux.scala 19:72:@31200.4]
  wire [7:0] _T_60989; // @[Mux.scala 19:72:@31207.4]
  wire [15:0] _T_60990; // @[Mux.scala 19:72:@31208.4]
  wire [15:0] _T_60992; // @[Mux.scala 19:72:@31209.4]
  wire [7:0] _T_60999; // @[Mux.scala 19:72:@31216.4]
  wire [7:0] _T_61006; // @[Mux.scala 19:72:@31223.4]
  wire [15:0] _T_61007; // @[Mux.scala 19:72:@31224.4]
  wire [15:0] _T_61009; // @[Mux.scala 19:72:@31225.4]
  wire [7:0] _T_61016; // @[Mux.scala 19:72:@31232.4]
  wire [7:0] _T_61023; // @[Mux.scala 19:72:@31239.4]
  wire [15:0] _T_61024; // @[Mux.scala 19:72:@31240.4]
  wire [15:0] _T_61026; // @[Mux.scala 19:72:@31241.4]
  wire [7:0] _T_61033; // @[Mux.scala 19:72:@31248.4]
  wire [7:0] _T_61040; // @[Mux.scala 19:72:@31255.4]
  wire [15:0] _T_61041; // @[Mux.scala 19:72:@31256.4]
  wire [15:0] _T_61043; // @[Mux.scala 19:72:@31257.4]
  wire [15:0] _T_61058; // @[Mux.scala 19:72:@31272.4]
  wire [15:0] _T_61060; // @[Mux.scala 19:72:@31273.4]
  wire [15:0] _T_61075; // @[Mux.scala 19:72:@31288.4]
  wire [15:0] _T_61077; // @[Mux.scala 19:72:@31289.4]
  wire [15:0] _T_61092; // @[Mux.scala 19:72:@31304.4]
  wire [15:0] _T_61094; // @[Mux.scala 19:72:@31305.4]
  wire [15:0] _T_61109; // @[Mux.scala 19:72:@31320.4]
  wire [15:0] _T_61111; // @[Mux.scala 19:72:@31321.4]
  wire [15:0] _T_61126; // @[Mux.scala 19:72:@31336.4]
  wire [15:0] _T_61128; // @[Mux.scala 19:72:@31337.4]
  wire [15:0] _T_61143; // @[Mux.scala 19:72:@31352.4]
  wire [15:0] _T_61145; // @[Mux.scala 19:72:@31353.4]
  wire [15:0] _T_61160; // @[Mux.scala 19:72:@31368.4]
  wire [15:0] _T_61162; // @[Mux.scala 19:72:@31369.4]
  wire [15:0] _T_61177; // @[Mux.scala 19:72:@31384.4]
  wire [15:0] _T_61179; // @[Mux.scala 19:72:@31385.4]
  wire [15:0] _T_61180; // @[Mux.scala 19:72:@31386.4]
  wire [15:0] _T_61181; // @[Mux.scala 19:72:@31387.4]
  wire [15:0] _T_61182; // @[Mux.scala 19:72:@31388.4]
  wire [15:0] _T_61183; // @[Mux.scala 19:72:@31389.4]
  wire [15:0] _T_61184; // @[Mux.scala 19:72:@31390.4]
  wire [15:0] _T_61185; // @[Mux.scala 19:72:@31391.4]
  wire [15:0] _T_61186; // @[Mux.scala 19:72:@31392.4]
  wire [15:0] _T_61187; // @[Mux.scala 19:72:@31393.4]
  wire [15:0] _T_61188; // @[Mux.scala 19:72:@31394.4]
  wire [15:0] _T_61189; // @[Mux.scala 19:72:@31395.4]
  wire [15:0] _T_61190; // @[Mux.scala 19:72:@31396.4]
  wire [15:0] _T_61191; // @[Mux.scala 19:72:@31397.4]
  wire [15:0] _T_61192; // @[Mux.scala 19:72:@31398.4]
  wire [15:0] _T_61193; // @[Mux.scala 19:72:@31399.4]
  wire [15:0] _T_61194; // @[Mux.scala 19:72:@31400.4]
  wire [7:0] _T_61772; // @[Mux.scala 19:72:@31750.4]
  wire [7:0] _T_61779; // @[Mux.scala 19:72:@31757.4]
  wire [15:0] _T_61780; // @[Mux.scala 19:72:@31758.4]
  wire [15:0] _T_61782; // @[Mux.scala 19:72:@31759.4]
  wire [7:0] _T_61789; // @[Mux.scala 19:72:@31766.4]
  wire [7:0] _T_61796; // @[Mux.scala 19:72:@31773.4]
  wire [15:0] _T_61797; // @[Mux.scala 19:72:@31774.4]
  wire [15:0] _T_61799; // @[Mux.scala 19:72:@31775.4]
  wire [7:0] _T_61806; // @[Mux.scala 19:72:@31782.4]
  wire [7:0] _T_61813; // @[Mux.scala 19:72:@31789.4]
  wire [15:0] _T_61814; // @[Mux.scala 19:72:@31790.4]
  wire [15:0] _T_61816; // @[Mux.scala 19:72:@31791.4]
  wire [7:0] _T_61823; // @[Mux.scala 19:72:@31798.4]
  wire [7:0] _T_61830; // @[Mux.scala 19:72:@31805.4]
  wire [15:0] _T_61831; // @[Mux.scala 19:72:@31806.4]
  wire [15:0] _T_61833; // @[Mux.scala 19:72:@31807.4]
  wire [7:0] _T_61840; // @[Mux.scala 19:72:@31814.4]
  wire [7:0] _T_61847; // @[Mux.scala 19:72:@31821.4]
  wire [15:0] _T_61848; // @[Mux.scala 19:72:@31822.4]
  wire [15:0] _T_61850; // @[Mux.scala 19:72:@31823.4]
  wire [7:0] _T_61857; // @[Mux.scala 19:72:@31830.4]
  wire [7:0] _T_61864; // @[Mux.scala 19:72:@31837.4]
  wire [15:0] _T_61865; // @[Mux.scala 19:72:@31838.4]
  wire [15:0] _T_61867; // @[Mux.scala 19:72:@31839.4]
  wire [7:0] _T_61874; // @[Mux.scala 19:72:@31846.4]
  wire [7:0] _T_61881; // @[Mux.scala 19:72:@31853.4]
  wire [15:0] _T_61882; // @[Mux.scala 19:72:@31854.4]
  wire [15:0] _T_61884; // @[Mux.scala 19:72:@31855.4]
  wire [7:0] _T_61891; // @[Mux.scala 19:72:@31862.4]
  wire [7:0] _T_61898; // @[Mux.scala 19:72:@31869.4]
  wire [15:0] _T_61899; // @[Mux.scala 19:72:@31870.4]
  wire [15:0] _T_61901; // @[Mux.scala 19:72:@31871.4]
  wire [15:0] _T_61916; // @[Mux.scala 19:72:@31886.4]
  wire [15:0] _T_61918; // @[Mux.scala 19:72:@31887.4]
  wire [15:0] _T_61933; // @[Mux.scala 19:72:@31902.4]
  wire [15:0] _T_61935; // @[Mux.scala 19:72:@31903.4]
  wire [15:0] _T_61950; // @[Mux.scala 19:72:@31918.4]
  wire [15:0] _T_61952; // @[Mux.scala 19:72:@31919.4]
  wire [15:0] _T_61967; // @[Mux.scala 19:72:@31934.4]
  wire [15:0] _T_61969; // @[Mux.scala 19:72:@31935.4]
  wire [15:0] _T_61984; // @[Mux.scala 19:72:@31950.4]
  wire [15:0] _T_61986; // @[Mux.scala 19:72:@31951.4]
  wire [15:0] _T_62001; // @[Mux.scala 19:72:@31966.4]
  wire [15:0] _T_62003; // @[Mux.scala 19:72:@31967.4]
  wire [15:0] _T_62018; // @[Mux.scala 19:72:@31982.4]
  wire [15:0] _T_62020; // @[Mux.scala 19:72:@31983.4]
  wire [15:0] _T_62035; // @[Mux.scala 19:72:@31998.4]
  wire [15:0] _T_62037; // @[Mux.scala 19:72:@31999.4]
  wire [15:0] _T_62038; // @[Mux.scala 19:72:@32000.4]
  wire [15:0] _T_62039; // @[Mux.scala 19:72:@32001.4]
  wire [15:0] _T_62040; // @[Mux.scala 19:72:@32002.4]
  wire [15:0] _T_62041; // @[Mux.scala 19:72:@32003.4]
  wire [15:0] _T_62042; // @[Mux.scala 19:72:@32004.4]
  wire [15:0] _T_62043; // @[Mux.scala 19:72:@32005.4]
  wire [15:0] _T_62044; // @[Mux.scala 19:72:@32006.4]
  wire [15:0] _T_62045; // @[Mux.scala 19:72:@32007.4]
  wire [15:0] _T_62046; // @[Mux.scala 19:72:@32008.4]
  wire [15:0] _T_62047; // @[Mux.scala 19:72:@32009.4]
  wire [15:0] _T_62048; // @[Mux.scala 19:72:@32010.4]
  wire [15:0] _T_62049; // @[Mux.scala 19:72:@32011.4]
  wire [15:0] _T_62050; // @[Mux.scala 19:72:@32012.4]
  wire [15:0] _T_62051; // @[Mux.scala 19:72:@32013.4]
  wire [15:0] _T_62052; // @[Mux.scala 19:72:@32014.4]
  wire [7:0] _T_62630; // @[Mux.scala 19:72:@32364.4]
  wire [7:0] _T_62637; // @[Mux.scala 19:72:@32371.4]
  wire [15:0] _T_62638; // @[Mux.scala 19:72:@32372.4]
  wire [15:0] _T_62640; // @[Mux.scala 19:72:@32373.4]
  wire [7:0] _T_62647; // @[Mux.scala 19:72:@32380.4]
  wire [7:0] _T_62654; // @[Mux.scala 19:72:@32387.4]
  wire [15:0] _T_62655; // @[Mux.scala 19:72:@32388.4]
  wire [15:0] _T_62657; // @[Mux.scala 19:72:@32389.4]
  wire [7:0] _T_62664; // @[Mux.scala 19:72:@32396.4]
  wire [7:0] _T_62671; // @[Mux.scala 19:72:@32403.4]
  wire [15:0] _T_62672; // @[Mux.scala 19:72:@32404.4]
  wire [15:0] _T_62674; // @[Mux.scala 19:72:@32405.4]
  wire [7:0] _T_62681; // @[Mux.scala 19:72:@32412.4]
  wire [7:0] _T_62688; // @[Mux.scala 19:72:@32419.4]
  wire [15:0] _T_62689; // @[Mux.scala 19:72:@32420.4]
  wire [15:0] _T_62691; // @[Mux.scala 19:72:@32421.4]
  wire [7:0] _T_62698; // @[Mux.scala 19:72:@32428.4]
  wire [7:0] _T_62705; // @[Mux.scala 19:72:@32435.4]
  wire [15:0] _T_62706; // @[Mux.scala 19:72:@32436.4]
  wire [15:0] _T_62708; // @[Mux.scala 19:72:@32437.4]
  wire [7:0] _T_62715; // @[Mux.scala 19:72:@32444.4]
  wire [7:0] _T_62722; // @[Mux.scala 19:72:@32451.4]
  wire [15:0] _T_62723; // @[Mux.scala 19:72:@32452.4]
  wire [15:0] _T_62725; // @[Mux.scala 19:72:@32453.4]
  wire [7:0] _T_62732; // @[Mux.scala 19:72:@32460.4]
  wire [7:0] _T_62739; // @[Mux.scala 19:72:@32467.4]
  wire [15:0] _T_62740; // @[Mux.scala 19:72:@32468.4]
  wire [15:0] _T_62742; // @[Mux.scala 19:72:@32469.4]
  wire [7:0] _T_62749; // @[Mux.scala 19:72:@32476.4]
  wire [7:0] _T_62756; // @[Mux.scala 19:72:@32483.4]
  wire [15:0] _T_62757; // @[Mux.scala 19:72:@32484.4]
  wire [15:0] _T_62759; // @[Mux.scala 19:72:@32485.4]
  wire [15:0] _T_62774; // @[Mux.scala 19:72:@32500.4]
  wire [15:0] _T_62776; // @[Mux.scala 19:72:@32501.4]
  wire [15:0] _T_62791; // @[Mux.scala 19:72:@32516.4]
  wire [15:0] _T_62793; // @[Mux.scala 19:72:@32517.4]
  wire [15:0] _T_62808; // @[Mux.scala 19:72:@32532.4]
  wire [15:0] _T_62810; // @[Mux.scala 19:72:@32533.4]
  wire [15:0] _T_62825; // @[Mux.scala 19:72:@32548.4]
  wire [15:0] _T_62827; // @[Mux.scala 19:72:@32549.4]
  wire [15:0] _T_62842; // @[Mux.scala 19:72:@32564.4]
  wire [15:0] _T_62844; // @[Mux.scala 19:72:@32565.4]
  wire [15:0] _T_62859; // @[Mux.scala 19:72:@32580.4]
  wire [15:0] _T_62861; // @[Mux.scala 19:72:@32581.4]
  wire [15:0] _T_62876; // @[Mux.scala 19:72:@32596.4]
  wire [15:0] _T_62878; // @[Mux.scala 19:72:@32597.4]
  wire [15:0] _T_62893; // @[Mux.scala 19:72:@32612.4]
  wire [15:0] _T_62895; // @[Mux.scala 19:72:@32613.4]
  wire [15:0] _T_62896; // @[Mux.scala 19:72:@32614.4]
  wire [15:0] _T_62897; // @[Mux.scala 19:72:@32615.4]
  wire [15:0] _T_62898; // @[Mux.scala 19:72:@32616.4]
  wire [15:0] _T_62899; // @[Mux.scala 19:72:@32617.4]
  wire [15:0] _T_62900; // @[Mux.scala 19:72:@32618.4]
  wire [15:0] _T_62901; // @[Mux.scala 19:72:@32619.4]
  wire [15:0] _T_62902; // @[Mux.scala 19:72:@32620.4]
  wire [15:0] _T_62903; // @[Mux.scala 19:72:@32621.4]
  wire [15:0] _T_62904; // @[Mux.scala 19:72:@32622.4]
  wire [15:0] _T_62905; // @[Mux.scala 19:72:@32623.4]
  wire [15:0] _T_62906; // @[Mux.scala 19:72:@32624.4]
  wire [15:0] _T_62907; // @[Mux.scala 19:72:@32625.4]
  wire [15:0] _T_62908; // @[Mux.scala 19:72:@32626.4]
  wire [15:0] _T_62909; // @[Mux.scala 19:72:@32627.4]
  wire [15:0] _T_62910; // @[Mux.scala 19:72:@32628.4]
  wire [7:0] _T_63488; // @[Mux.scala 19:72:@32978.4]
  wire [7:0] _T_63495; // @[Mux.scala 19:72:@32985.4]
  wire [15:0] _T_63496; // @[Mux.scala 19:72:@32986.4]
  wire [15:0] _T_63498; // @[Mux.scala 19:72:@32987.4]
  wire [7:0] _T_63505; // @[Mux.scala 19:72:@32994.4]
  wire [7:0] _T_63512; // @[Mux.scala 19:72:@33001.4]
  wire [15:0] _T_63513; // @[Mux.scala 19:72:@33002.4]
  wire [15:0] _T_63515; // @[Mux.scala 19:72:@33003.4]
  wire [7:0] _T_63522; // @[Mux.scala 19:72:@33010.4]
  wire [7:0] _T_63529; // @[Mux.scala 19:72:@33017.4]
  wire [15:0] _T_63530; // @[Mux.scala 19:72:@33018.4]
  wire [15:0] _T_63532; // @[Mux.scala 19:72:@33019.4]
  wire [7:0] _T_63539; // @[Mux.scala 19:72:@33026.4]
  wire [7:0] _T_63546; // @[Mux.scala 19:72:@33033.4]
  wire [15:0] _T_63547; // @[Mux.scala 19:72:@33034.4]
  wire [15:0] _T_63549; // @[Mux.scala 19:72:@33035.4]
  wire [7:0] _T_63556; // @[Mux.scala 19:72:@33042.4]
  wire [7:0] _T_63563; // @[Mux.scala 19:72:@33049.4]
  wire [15:0] _T_63564; // @[Mux.scala 19:72:@33050.4]
  wire [15:0] _T_63566; // @[Mux.scala 19:72:@33051.4]
  wire [7:0] _T_63573; // @[Mux.scala 19:72:@33058.4]
  wire [7:0] _T_63580; // @[Mux.scala 19:72:@33065.4]
  wire [15:0] _T_63581; // @[Mux.scala 19:72:@33066.4]
  wire [15:0] _T_63583; // @[Mux.scala 19:72:@33067.4]
  wire [7:0] _T_63590; // @[Mux.scala 19:72:@33074.4]
  wire [7:0] _T_63597; // @[Mux.scala 19:72:@33081.4]
  wire [15:0] _T_63598; // @[Mux.scala 19:72:@33082.4]
  wire [15:0] _T_63600; // @[Mux.scala 19:72:@33083.4]
  wire [7:0] _T_63607; // @[Mux.scala 19:72:@33090.4]
  wire [7:0] _T_63614; // @[Mux.scala 19:72:@33097.4]
  wire [15:0] _T_63615; // @[Mux.scala 19:72:@33098.4]
  wire [15:0] _T_63617; // @[Mux.scala 19:72:@33099.4]
  wire [15:0] _T_63632; // @[Mux.scala 19:72:@33114.4]
  wire [15:0] _T_63634; // @[Mux.scala 19:72:@33115.4]
  wire [15:0] _T_63649; // @[Mux.scala 19:72:@33130.4]
  wire [15:0] _T_63651; // @[Mux.scala 19:72:@33131.4]
  wire [15:0] _T_63666; // @[Mux.scala 19:72:@33146.4]
  wire [15:0] _T_63668; // @[Mux.scala 19:72:@33147.4]
  wire [15:0] _T_63683; // @[Mux.scala 19:72:@33162.4]
  wire [15:0] _T_63685; // @[Mux.scala 19:72:@33163.4]
  wire [15:0] _T_63700; // @[Mux.scala 19:72:@33178.4]
  wire [15:0] _T_63702; // @[Mux.scala 19:72:@33179.4]
  wire [15:0] _T_63717; // @[Mux.scala 19:72:@33194.4]
  wire [15:0] _T_63719; // @[Mux.scala 19:72:@33195.4]
  wire [15:0] _T_63734; // @[Mux.scala 19:72:@33210.4]
  wire [15:0] _T_63736; // @[Mux.scala 19:72:@33211.4]
  wire [15:0] _T_63751; // @[Mux.scala 19:72:@33226.4]
  wire [15:0] _T_63753; // @[Mux.scala 19:72:@33227.4]
  wire [15:0] _T_63754; // @[Mux.scala 19:72:@33228.4]
  wire [15:0] _T_63755; // @[Mux.scala 19:72:@33229.4]
  wire [15:0] _T_63756; // @[Mux.scala 19:72:@33230.4]
  wire [15:0] _T_63757; // @[Mux.scala 19:72:@33231.4]
  wire [15:0] _T_63758; // @[Mux.scala 19:72:@33232.4]
  wire [15:0] _T_63759; // @[Mux.scala 19:72:@33233.4]
  wire [15:0] _T_63760; // @[Mux.scala 19:72:@33234.4]
  wire [15:0] _T_63761; // @[Mux.scala 19:72:@33235.4]
  wire [15:0] _T_63762; // @[Mux.scala 19:72:@33236.4]
  wire [15:0] _T_63763; // @[Mux.scala 19:72:@33237.4]
  wire [15:0] _T_63764; // @[Mux.scala 19:72:@33238.4]
  wire [15:0] _T_63765; // @[Mux.scala 19:72:@33239.4]
  wire [15:0] _T_63766; // @[Mux.scala 19:72:@33240.4]
  wire [15:0] _T_63767; // @[Mux.scala 19:72:@33241.4]
  wire [15:0] _T_63768; // @[Mux.scala 19:72:@33242.4]
  wire [7:0] _T_64346; // @[Mux.scala 19:72:@33592.4]
  wire [7:0] _T_64353; // @[Mux.scala 19:72:@33599.4]
  wire [15:0] _T_64354; // @[Mux.scala 19:72:@33600.4]
  wire [15:0] _T_64356; // @[Mux.scala 19:72:@33601.4]
  wire [7:0] _T_64363; // @[Mux.scala 19:72:@33608.4]
  wire [7:0] _T_64370; // @[Mux.scala 19:72:@33615.4]
  wire [15:0] _T_64371; // @[Mux.scala 19:72:@33616.4]
  wire [15:0] _T_64373; // @[Mux.scala 19:72:@33617.4]
  wire [7:0] _T_64380; // @[Mux.scala 19:72:@33624.4]
  wire [7:0] _T_64387; // @[Mux.scala 19:72:@33631.4]
  wire [15:0] _T_64388; // @[Mux.scala 19:72:@33632.4]
  wire [15:0] _T_64390; // @[Mux.scala 19:72:@33633.4]
  wire [7:0] _T_64397; // @[Mux.scala 19:72:@33640.4]
  wire [7:0] _T_64404; // @[Mux.scala 19:72:@33647.4]
  wire [15:0] _T_64405; // @[Mux.scala 19:72:@33648.4]
  wire [15:0] _T_64407; // @[Mux.scala 19:72:@33649.4]
  wire [7:0] _T_64414; // @[Mux.scala 19:72:@33656.4]
  wire [7:0] _T_64421; // @[Mux.scala 19:72:@33663.4]
  wire [15:0] _T_64422; // @[Mux.scala 19:72:@33664.4]
  wire [15:0] _T_64424; // @[Mux.scala 19:72:@33665.4]
  wire [7:0] _T_64431; // @[Mux.scala 19:72:@33672.4]
  wire [7:0] _T_64438; // @[Mux.scala 19:72:@33679.4]
  wire [15:0] _T_64439; // @[Mux.scala 19:72:@33680.4]
  wire [15:0] _T_64441; // @[Mux.scala 19:72:@33681.4]
  wire [7:0] _T_64448; // @[Mux.scala 19:72:@33688.4]
  wire [7:0] _T_64455; // @[Mux.scala 19:72:@33695.4]
  wire [15:0] _T_64456; // @[Mux.scala 19:72:@33696.4]
  wire [15:0] _T_64458; // @[Mux.scala 19:72:@33697.4]
  wire [7:0] _T_64465; // @[Mux.scala 19:72:@33704.4]
  wire [7:0] _T_64472; // @[Mux.scala 19:72:@33711.4]
  wire [15:0] _T_64473; // @[Mux.scala 19:72:@33712.4]
  wire [15:0] _T_64475; // @[Mux.scala 19:72:@33713.4]
  wire [15:0] _T_64490; // @[Mux.scala 19:72:@33728.4]
  wire [15:0] _T_64492; // @[Mux.scala 19:72:@33729.4]
  wire [15:0] _T_64507; // @[Mux.scala 19:72:@33744.4]
  wire [15:0] _T_64509; // @[Mux.scala 19:72:@33745.4]
  wire [15:0] _T_64524; // @[Mux.scala 19:72:@33760.4]
  wire [15:0] _T_64526; // @[Mux.scala 19:72:@33761.4]
  wire [15:0] _T_64541; // @[Mux.scala 19:72:@33776.4]
  wire [15:0] _T_64543; // @[Mux.scala 19:72:@33777.4]
  wire [15:0] _T_64558; // @[Mux.scala 19:72:@33792.4]
  wire [15:0] _T_64560; // @[Mux.scala 19:72:@33793.4]
  wire [15:0] _T_64575; // @[Mux.scala 19:72:@33808.4]
  wire [15:0] _T_64577; // @[Mux.scala 19:72:@33809.4]
  wire [15:0] _T_64592; // @[Mux.scala 19:72:@33824.4]
  wire [15:0] _T_64594; // @[Mux.scala 19:72:@33825.4]
  wire [15:0] _T_64609; // @[Mux.scala 19:72:@33840.4]
  wire [15:0] _T_64611; // @[Mux.scala 19:72:@33841.4]
  wire [15:0] _T_64612; // @[Mux.scala 19:72:@33842.4]
  wire [15:0] _T_64613; // @[Mux.scala 19:72:@33843.4]
  wire [15:0] _T_64614; // @[Mux.scala 19:72:@33844.4]
  wire [15:0] _T_64615; // @[Mux.scala 19:72:@33845.4]
  wire [15:0] _T_64616; // @[Mux.scala 19:72:@33846.4]
  wire [15:0] _T_64617; // @[Mux.scala 19:72:@33847.4]
  wire [15:0] _T_64618; // @[Mux.scala 19:72:@33848.4]
  wire [15:0] _T_64619; // @[Mux.scala 19:72:@33849.4]
  wire [15:0] _T_64620; // @[Mux.scala 19:72:@33850.4]
  wire [15:0] _T_64621; // @[Mux.scala 19:72:@33851.4]
  wire [15:0] _T_64622; // @[Mux.scala 19:72:@33852.4]
  wire [15:0] _T_64623; // @[Mux.scala 19:72:@33853.4]
  wire [15:0] _T_64624; // @[Mux.scala 19:72:@33854.4]
  wire [15:0] _T_64625; // @[Mux.scala 19:72:@33855.4]
  wire [15:0] _T_64626; // @[Mux.scala 19:72:@33856.4]
  wire [7:0] _T_65204; // @[Mux.scala 19:72:@34206.4]
  wire [7:0] _T_65211; // @[Mux.scala 19:72:@34213.4]
  wire [15:0] _T_65212; // @[Mux.scala 19:72:@34214.4]
  wire [15:0] _T_65214; // @[Mux.scala 19:72:@34215.4]
  wire [7:0] _T_65221; // @[Mux.scala 19:72:@34222.4]
  wire [7:0] _T_65228; // @[Mux.scala 19:72:@34229.4]
  wire [15:0] _T_65229; // @[Mux.scala 19:72:@34230.4]
  wire [15:0] _T_65231; // @[Mux.scala 19:72:@34231.4]
  wire [7:0] _T_65238; // @[Mux.scala 19:72:@34238.4]
  wire [7:0] _T_65245; // @[Mux.scala 19:72:@34245.4]
  wire [15:0] _T_65246; // @[Mux.scala 19:72:@34246.4]
  wire [15:0] _T_65248; // @[Mux.scala 19:72:@34247.4]
  wire [7:0] _T_65255; // @[Mux.scala 19:72:@34254.4]
  wire [7:0] _T_65262; // @[Mux.scala 19:72:@34261.4]
  wire [15:0] _T_65263; // @[Mux.scala 19:72:@34262.4]
  wire [15:0] _T_65265; // @[Mux.scala 19:72:@34263.4]
  wire [7:0] _T_65272; // @[Mux.scala 19:72:@34270.4]
  wire [7:0] _T_65279; // @[Mux.scala 19:72:@34277.4]
  wire [15:0] _T_65280; // @[Mux.scala 19:72:@34278.4]
  wire [15:0] _T_65282; // @[Mux.scala 19:72:@34279.4]
  wire [7:0] _T_65289; // @[Mux.scala 19:72:@34286.4]
  wire [7:0] _T_65296; // @[Mux.scala 19:72:@34293.4]
  wire [15:0] _T_65297; // @[Mux.scala 19:72:@34294.4]
  wire [15:0] _T_65299; // @[Mux.scala 19:72:@34295.4]
  wire [7:0] _T_65306; // @[Mux.scala 19:72:@34302.4]
  wire [7:0] _T_65313; // @[Mux.scala 19:72:@34309.4]
  wire [15:0] _T_65314; // @[Mux.scala 19:72:@34310.4]
  wire [15:0] _T_65316; // @[Mux.scala 19:72:@34311.4]
  wire [7:0] _T_65323; // @[Mux.scala 19:72:@34318.4]
  wire [7:0] _T_65330; // @[Mux.scala 19:72:@34325.4]
  wire [15:0] _T_65331; // @[Mux.scala 19:72:@34326.4]
  wire [15:0] _T_65333; // @[Mux.scala 19:72:@34327.4]
  wire [15:0] _T_65348; // @[Mux.scala 19:72:@34342.4]
  wire [15:0] _T_65350; // @[Mux.scala 19:72:@34343.4]
  wire [15:0] _T_65365; // @[Mux.scala 19:72:@34358.4]
  wire [15:0] _T_65367; // @[Mux.scala 19:72:@34359.4]
  wire [15:0] _T_65382; // @[Mux.scala 19:72:@34374.4]
  wire [15:0] _T_65384; // @[Mux.scala 19:72:@34375.4]
  wire [15:0] _T_65399; // @[Mux.scala 19:72:@34390.4]
  wire [15:0] _T_65401; // @[Mux.scala 19:72:@34391.4]
  wire [15:0] _T_65416; // @[Mux.scala 19:72:@34406.4]
  wire [15:0] _T_65418; // @[Mux.scala 19:72:@34407.4]
  wire [15:0] _T_65433; // @[Mux.scala 19:72:@34422.4]
  wire [15:0] _T_65435; // @[Mux.scala 19:72:@34423.4]
  wire [15:0] _T_65450; // @[Mux.scala 19:72:@34438.4]
  wire [15:0] _T_65452; // @[Mux.scala 19:72:@34439.4]
  wire [15:0] _T_65467; // @[Mux.scala 19:72:@34454.4]
  wire [15:0] _T_65469; // @[Mux.scala 19:72:@34455.4]
  wire [15:0] _T_65470; // @[Mux.scala 19:72:@34456.4]
  wire [15:0] _T_65471; // @[Mux.scala 19:72:@34457.4]
  wire [15:0] _T_65472; // @[Mux.scala 19:72:@34458.4]
  wire [15:0] _T_65473; // @[Mux.scala 19:72:@34459.4]
  wire [15:0] _T_65474; // @[Mux.scala 19:72:@34460.4]
  wire [15:0] _T_65475; // @[Mux.scala 19:72:@34461.4]
  wire [15:0] _T_65476; // @[Mux.scala 19:72:@34462.4]
  wire [15:0] _T_65477; // @[Mux.scala 19:72:@34463.4]
  wire [15:0] _T_65478; // @[Mux.scala 19:72:@34464.4]
  wire [15:0] _T_65479; // @[Mux.scala 19:72:@34465.4]
  wire [15:0] _T_65480; // @[Mux.scala 19:72:@34466.4]
  wire [15:0] _T_65481; // @[Mux.scala 19:72:@34467.4]
  wire [15:0] _T_65482; // @[Mux.scala 19:72:@34468.4]
  wire [15:0] _T_65483; // @[Mux.scala 19:72:@34469.4]
  wire [15:0] _T_65484; // @[Mux.scala 19:72:@34470.4]
  reg  storeAddrNotKnownFlagsPReg_0_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_419;
  reg  storeAddrNotKnownFlagsPReg_0_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_420;
  reg  storeAddrNotKnownFlagsPReg_0_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_421;
  reg  storeAddrNotKnownFlagsPReg_0_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_422;
  reg  storeAddrNotKnownFlagsPReg_0_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_423;
  reg  storeAddrNotKnownFlagsPReg_0_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_424;
  reg  storeAddrNotKnownFlagsPReg_0_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_425;
  reg  storeAddrNotKnownFlagsPReg_0_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_426;
  reg  storeAddrNotKnownFlagsPReg_0_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_427;
  reg  storeAddrNotKnownFlagsPReg_0_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_428;
  reg  storeAddrNotKnownFlagsPReg_0_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_429;
  reg  storeAddrNotKnownFlagsPReg_0_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_430;
  reg  storeAddrNotKnownFlagsPReg_0_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_431;
  reg  storeAddrNotKnownFlagsPReg_0_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_432;
  reg  storeAddrNotKnownFlagsPReg_0_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_433;
  reg  storeAddrNotKnownFlagsPReg_0_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_434;
  reg  storeAddrNotKnownFlagsPReg_1_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_435;
  reg  storeAddrNotKnownFlagsPReg_1_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_436;
  reg  storeAddrNotKnownFlagsPReg_1_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_437;
  reg  storeAddrNotKnownFlagsPReg_1_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_438;
  reg  storeAddrNotKnownFlagsPReg_1_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_439;
  reg  storeAddrNotKnownFlagsPReg_1_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_440;
  reg  storeAddrNotKnownFlagsPReg_1_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_441;
  reg  storeAddrNotKnownFlagsPReg_1_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_442;
  reg  storeAddrNotKnownFlagsPReg_1_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_443;
  reg  storeAddrNotKnownFlagsPReg_1_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_444;
  reg  storeAddrNotKnownFlagsPReg_1_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_445;
  reg  storeAddrNotKnownFlagsPReg_1_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_446;
  reg  storeAddrNotKnownFlagsPReg_1_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_447;
  reg  storeAddrNotKnownFlagsPReg_1_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_448;
  reg  storeAddrNotKnownFlagsPReg_1_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_449;
  reg  storeAddrNotKnownFlagsPReg_1_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_450;
  reg  storeAddrNotKnownFlagsPReg_2_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_451;
  reg  storeAddrNotKnownFlagsPReg_2_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_452;
  reg  storeAddrNotKnownFlagsPReg_2_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_453;
  reg  storeAddrNotKnownFlagsPReg_2_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_454;
  reg  storeAddrNotKnownFlagsPReg_2_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_455;
  reg  storeAddrNotKnownFlagsPReg_2_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_456;
  reg  storeAddrNotKnownFlagsPReg_2_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_457;
  reg  storeAddrNotKnownFlagsPReg_2_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_458;
  reg  storeAddrNotKnownFlagsPReg_2_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_459;
  reg  storeAddrNotKnownFlagsPReg_2_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_460;
  reg  storeAddrNotKnownFlagsPReg_2_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_461;
  reg  storeAddrNotKnownFlagsPReg_2_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_462;
  reg  storeAddrNotKnownFlagsPReg_2_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_463;
  reg  storeAddrNotKnownFlagsPReg_2_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_464;
  reg  storeAddrNotKnownFlagsPReg_2_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_465;
  reg  storeAddrNotKnownFlagsPReg_2_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_466;
  reg  storeAddrNotKnownFlagsPReg_3_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_467;
  reg  storeAddrNotKnownFlagsPReg_3_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_468;
  reg  storeAddrNotKnownFlagsPReg_3_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_469;
  reg  storeAddrNotKnownFlagsPReg_3_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_470;
  reg  storeAddrNotKnownFlagsPReg_3_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_471;
  reg  storeAddrNotKnownFlagsPReg_3_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_472;
  reg  storeAddrNotKnownFlagsPReg_3_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_473;
  reg  storeAddrNotKnownFlagsPReg_3_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_474;
  reg  storeAddrNotKnownFlagsPReg_3_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_475;
  reg  storeAddrNotKnownFlagsPReg_3_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_476;
  reg  storeAddrNotKnownFlagsPReg_3_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_477;
  reg  storeAddrNotKnownFlagsPReg_3_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_478;
  reg  storeAddrNotKnownFlagsPReg_3_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_479;
  reg  storeAddrNotKnownFlagsPReg_3_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_480;
  reg  storeAddrNotKnownFlagsPReg_3_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_481;
  reg  storeAddrNotKnownFlagsPReg_3_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_482;
  reg  storeAddrNotKnownFlagsPReg_4_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_483;
  reg  storeAddrNotKnownFlagsPReg_4_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_484;
  reg  storeAddrNotKnownFlagsPReg_4_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_485;
  reg  storeAddrNotKnownFlagsPReg_4_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_486;
  reg  storeAddrNotKnownFlagsPReg_4_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_487;
  reg  storeAddrNotKnownFlagsPReg_4_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_488;
  reg  storeAddrNotKnownFlagsPReg_4_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_489;
  reg  storeAddrNotKnownFlagsPReg_4_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_490;
  reg  storeAddrNotKnownFlagsPReg_4_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_491;
  reg  storeAddrNotKnownFlagsPReg_4_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_492;
  reg  storeAddrNotKnownFlagsPReg_4_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_493;
  reg  storeAddrNotKnownFlagsPReg_4_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_494;
  reg  storeAddrNotKnownFlagsPReg_4_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_495;
  reg  storeAddrNotKnownFlagsPReg_4_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_496;
  reg  storeAddrNotKnownFlagsPReg_4_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_497;
  reg  storeAddrNotKnownFlagsPReg_4_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_498;
  reg  storeAddrNotKnownFlagsPReg_5_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_499;
  reg  storeAddrNotKnownFlagsPReg_5_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_500;
  reg  storeAddrNotKnownFlagsPReg_5_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_501;
  reg  storeAddrNotKnownFlagsPReg_5_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_502;
  reg  storeAddrNotKnownFlagsPReg_5_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_503;
  reg  storeAddrNotKnownFlagsPReg_5_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_504;
  reg  storeAddrNotKnownFlagsPReg_5_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_505;
  reg  storeAddrNotKnownFlagsPReg_5_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_506;
  reg  storeAddrNotKnownFlagsPReg_5_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_507;
  reg  storeAddrNotKnownFlagsPReg_5_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_508;
  reg  storeAddrNotKnownFlagsPReg_5_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_509;
  reg  storeAddrNotKnownFlagsPReg_5_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_510;
  reg  storeAddrNotKnownFlagsPReg_5_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_511;
  reg  storeAddrNotKnownFlagsPReg_5_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_512;
  reg  storeAddrNotKnownFlagsPReg_5_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_513;
  reg  storeAddrNotKnownFlagsPReg_5_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_514;
  reg  storeAddrNotKnownFlagsPReg_6_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_515;
  reg  storeAddrNotKnownFlagsPReg_6_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_516;
  reg  storeAddrNotKnownFlagsPReg_6_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_517;
  reg  storeAddrNotKnownFlagsPReg_6_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_518;
  reg  storeAddrNotKnownFlagsPReg_6_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_519;
  reg  storeAddrNotKnownFlagsPReg_6_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_520;
  reg  storeAddrNotKnownFlagsPReg_6_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_521;
  reg  storeAddrNotKnownFlagsPReg_6_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_522;
  reg  storeAddrNotKnownFlagsPReg_6_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_523;
  reg  storeAddrNotKnownFlagsPReg_6_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_524;
  reg  storeAddrNotKnownFlagsPReg_6_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_525;
  reg  storeAddrNotKnownFlagsPReg_6_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_526;
  reg  storeAddrNotKnownFlagsPReg_6_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_527;
  reg  storeAddrNotKnownFlagsPReg_6_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_528;
  reg  storeAddrNotKnownFlagsPReg_6_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_529;
  reg  storeAddrNotKnownFlagsPReg_6_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_530;
  reg  storeAddrNotKnownFlagsPReg_7_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_531;
  reg  storeAddrNotKnownFlagsPReg_7_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_532;
  reg  storeAddrNotKnownFlagsPReg_7_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_533;
  reg  storeAddrNotKnownFlagsPReg_7_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_534;
  reg  storeAddrNotKnownFlagsPReg_7_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_535;
  reg  storeAddrNotKnownFlagsPReg_7_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_536;
  reg  storeAddrNotKnownFlagsPReg_7_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_537;
  reg  storeAddrNotKnownFlagsPReg_7_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_538;
  reg  storeAddrNotKnownFlagsPReg_7_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_539;
  reg  storeAddrNotKnownFlagsPReg_7_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_540;
  reg  storeAddrNotKnownFlagsPReg_7_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_541;
  reg  storeAddrNotKnownFlagsPReg_7_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_542;
  reg  storeAddrNotKnownFlagsPReg_7_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_543;
  reg  storeAddrNotKnownFlagsPReg_7_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_544;
  reg  storeAddrNotKnownFlagsPReg_7_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_545;
  reg  storeAddrNotKnownFlagsPReg_7_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_546;
  reg  storeAddrNotKnownFlagsPReg_8_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_547;
  reg  storeAddrNotKnownFlagsPReg_8_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_548;
  reg  storeAddrNotKnownFlagsPReg_8_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_549;
  reg  storeAddrNotKnownFlagsPReg_8_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_550;
  reg  storeAddrNotKnownFlagsPReg_8_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_551;
  reg  storeAddrNotKnownFlagsPReg_8_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_552;
  reg  storeAddrNotKnownFlagsPReg_8_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_553;
  reg  storeAddrNotKnownFlagsPReg_8_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_554;
  reg  storeAddrNotKnownFlagsPReg_8_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_555;
  reg  storeAddrNotKnownFlagsPReg_8_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_556;
  reg  storeAddrNotKnownFlagsPReg_8_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_557;
  reg  storeAddrNotKnownFlagsPReg_8_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_558;
  reg  storeAddrNotKnownFlagsPReg_8_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_559;
  reg  storeAddrNotKnownFlagsPReg_8_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_560;
  reg  storeAddrNotKnownFlagsPReg_8_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_561;
  reg  storeAddrNotKnownFlagsPReg_8_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_562;
  reg  storeAddrNotKnownFlagsPReg_9_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_563;
  reg  storeAddrNotKnownFlagsPReg_9_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_564;
  reg  storeAddrNotKnownFlagsPReg_9_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_565;
  reg  storeAddrNotKnownFlagsPReg_9_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_566;
  reg  storeAddrNotKnownFlagsPReg_9_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_567;
  reg  storeAddrNotKnownFlagsPReg_9_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_568;
  reg  storeAddrNotKnownFlagsPReg_9_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_569;
  reg  storeAddrNotKnownFlagsPReg_9_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_570;
  reg  storeAddrNotKnownFlagsPReg_9_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_571;
  reg  storeAddrNotKnownFlagsPReg_9_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_572;
  reg  storeAddrNotKnownFlagsPReg_9_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_573;
  reg  storeAddrNotKnownFlagsPReg_9_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_574;
  reg  storeAddrNotKnownFlagsPReg_9_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_575;
  reg  storeAddrNotKnownFlagsPReg_9_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_576;
  reg  storeAddrNotKnownFlagsPReg_9_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_577;
  reg  storeAddrNotKnownFlagsPReg_9_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_578;
  reg  storeAddrNotKnownFlagsPReg_10_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_579;
  reg  storeAddrNotKnownFlagsPReg_10_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_580;
  reg  storeAddrNotKnownFlagsPReg_10_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_581;
  reg  storeAddrNotKnownFlagsPReg_10_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_582;
  reg  storeAddrNotKnownFlagsPReg_10_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_583;
  reg  storeAddrNotKnownFlagsPReg_10_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_584;
  reg  storeAddrNotKnownFlagsPReg_10_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_585;
  reg  storeAddrNotKnownFlagsPReg_10_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_586;
  reg  storeAddrNotKnownFlagsPReg_10_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_587;
  reg  storeAddrNotKnownFlagsPReg_10_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_588;
  reg  storeAddrNotKnownFlagsPReg_10_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_589;
  reg  storeAddrNotKnownFlagsPReg_10_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_590;
  reg  storeAddrNotKnownFlagsPReg_10_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_591;
  reg  storeAddrNotKnownFlagsPReg_10_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_592;
  reg  storeAddrNotKnownFlagsPReg_10_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_593;
  reg  storeAddrNotKnownFlagsPReg_10_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_594;
  reg  storeAddrNotKnownFlagsPReg_11_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_595;
  reg  storeAddrNotKnownFlagsPReg_11_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_596;
  reg  storeAddrNotKnownFlagsPReg_11_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_597;
  reg  storeAddrNotKnownFlagsPReg_11_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_598;
  reg  storeAddrNotKnownFlagsPReg_11_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_599;
  reg  storeAddrNotKnownFlagsPReg_11_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_600;
  reg  storeAddrNotKnownFlagsPReg_11_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_601;
  reg  storeAddrNotKnownFlagsPReg_11_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_602;
  reg  storeAddrNotKnownFlagsPReg_11_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_603;
  reg  storeAddrNotKnownFlagsPReg_11_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_604;
  reg  storeAddrNotKnownFlagsPReg_11_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_605;
  reg  storeAddrNotKnownFlagsPReg_11_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_606;
  reg  storeAddrNotKnownFlagsPReg_11_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_607;
  reg  storeAddrNotKnownFlagsPReg_11_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_608;
  reg  storeAddrNotKnownFlagsPReg_11_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_609;
  reg  storeAddrNotKnownFlagsPReg_11_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_610;
  reg  storeAddrNotKnownFlagsPReg_12_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_611;
  reg  storeAddrNotKnownFlagsPReg_12_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_612;
  reg  storeAddrNotKnownFlagsPReg_12_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_613;
  reg  storeAddrNotKnownFlagsPReg_12_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_614;
  reg  storeAddrNotKnownFlagsPReg_12_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_615;
  reg  storeAddrNotKnownFlagsPReg_12_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_616;
  reg  storeAddrNotKnownFlagsPReg_12_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_617;
  reg  storeAddrNotKnownFlagsPReg_12_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_618;
  reg  storeAddrNotKnownFlagsPReg_12_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_619;
  reg  storeAddrNotKnownFlagsPReg_12_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_620;
  reg  storeAddrNotKnownFlagsPReg_12_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_621;
  reg  storeAddrNotKnownFlagsPReg_12_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_622;
  reg  storeAddrNotKnownFlagsPReg_12_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_623;
  reg  storeAddrNotKnownFlagsPReg_12_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_624;
  reg  storeAddrNotKnownFlagsPReg_12_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_625;
  reg  storeAddrNotKnownFlagsPReg_12_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_626;
  reg  storeAddrNotKnownFlagsPReg_13_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_627;
  reg  storeAddrNotKnownFlagsPReg_13_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_628;
  reg  storeAddrNotKnownFlagsPReg_13_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_629;
  reg  storeAddrNotKnownFlagsPReg_13_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_630;
  reg  storeAddrNotKnownFlagsPReg_13_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_631;
  reg  storeAddrNotKnownFlagsPReg_13_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_632;
  reg  storeAddrNotKnownFlagsPReg_13_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_633;
  reg  storeAddrNotKnownFlagsPReg_13_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_634;
  reg  storeAddrNotKnownFlagsPReg_13_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_635;
  reg  storeAddrNotKnownFlagsPReg_13_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_636;
  reg  storeAddrNotKnownFlagsPReg_13_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_637;
  reg  storeAddrNotKnownFlagsPReg_13_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_638;
  reg  storeAddrNotKnownFlagsPReg_13_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_639;
  reg  storeAddrNotKnownFlagsPReg_13_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_640;
  reg  storeAddrNotKnownFlagsPReg_13_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_641;
  reg  storeAddrNotKnownFlagsPReg_13_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_642;
  reg  storeAddrNotKnownFlagsPReg_14_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_643;
  reg  storeAddrNotKnownFlagsPReg_14_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_644;
  reg  storeAddrNotKnownFlagsPReg_14_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_645;
  reg  storeAddrNotKnownFlagsPReg_14_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_646;
  reg  storeAddrNotKnownFlagsPReg_14_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_647;
  reg  storeAddrNotKnownFlagsPReg_14_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_648;
  reg  storeAddrNotKnownFlagsPReg_14_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_649;
  reg  storeAddrNotKnownFlagsPReg_14_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_650;
  reg  storeAddrNotKnownFlagsPReg_14_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_651;
  reg  storeAddrNotKnownFlagsPReg_14_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_652;
  reg  storeAddrNotKnownFlagsPReg_14_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_653;
  reg  storeAddrNotKnownFlagsPReg_14_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_654;
  reg  storeAddrNotKnownFlagsPReg_14_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_655;
  reg  storeAddrNotKnownFlagsPReg_14_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_656;
  reg  storeAddrNotKnownFlagsPReg_14_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_657;
  reg  storeAddrNotKnownFlagsPReg_14_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_658;
  reg  storeAddrNotKnownFlagsPReg_15_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_659;
  reg  storeAddrNotKnownFlagsPReg_15_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_660;
  reg  storeAddrNotKnownFlagsPReg_15_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_661;
  reg  storeAddrNotKnownFlagsPReg_15_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_662;
  reg  storeAddrNotKnownFlagsPReg_15_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_663;
  reg  storeAddrNotKnownFlagsPReg_15_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_664;
  reg  storeAddrNotKnownFlagsPReg_15_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_665;
  reg  storeAddrNotKnownFlagsPReg_15_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_666;
  reg  storeAddrNotKnownFlagsPReg_15_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_667;
  reg  storeAddrNotKnownFlagsPReg_15_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_668;
  reg  storeAddrNotKnownFlagsPReg_15_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_669;
  reg  storeAddrNotKnownFlagsPReg_15_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_670;
  reg  storeAddrNotKnownFlagsPReg_15_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_671;
  reg  storeAddrNotKnownFlagsPReg_15_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_672;
  reg  storeAddrNotKnownFlagsPReg_15_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_673;
  reg  storeAddrNotKnownFlagsPReg_15_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_674;
  reg  shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_675;
  reg  shiftedStoreDataKnownPReg_1; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_676;
  reg  shiftedStoreDataKnownPReg_2; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_677;
  reg  shiftedStoreDataKnownPReg_3; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_678;
  reg  shiftedStoreDataKnownPReg_4; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_679;
  reg  shiftedStoreDataKnownPReg_5; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_680;
  reg  shiftedStoreDataKnownPReg_6; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_681;
  reg  shiftedStoreDataKnownPReg_7; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_682;
  reg  shiftedStoreDataKnownPReg_8; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_683;
  reg  shiftedStoreDataKnownPReg_9; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_684;
  reg  shiftedStoreDataKnownPReg_10; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_685;
  reg  shiftedStoreDataKnownPReg_11; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_686;
  reg  shiftedStoreDataKnownPReg_12; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_687;
  reg  shiftedStoreDataKnownPReg_13; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_688;
  reg  shiftedStoreDataKnownPReg_14; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_689;
  reg  shiftedStoreDataKnownPReg_15; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_690;
  reg [31:0] shiftedStoreDataQPreg_0; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_691;
  reg [31:0] shiftedStoreDataQPreg_1; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_692;
  reg [31:0] shiftedStoreDataQPreg_2; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_693;
  reg [31:0] shiftedStoreDataQPreg_3; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_694;
  reg [31:0] shiftedStoreDataQPreg_4; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_695;
  reg [31:0] shiftedStoreDataQPreg_5; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_696;
  reg [31:0] shiftedStoreDataQPreg_6; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_697;
  reg [31:0] shiftedStoreDataQPreg_7; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_698;
  reg [31:0] shiftedStoreDataQPreg_8; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_699;
  reg [31:0] shiftedStoreDataQPreg_9; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_700;
  reg [31:0] shiftedStoreDataQPreg_10; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_701;
  reg [31:0] shiftedStoreDataQPreg_11; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_702;
  reg [31:0] shiftedStoreDataQPreg_12; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_703;
  reg [31:0] shiftedStoreDataQPreg_13; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_704;
  reg [31:0] shiftedStoreDataQPreg_14; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_705;
  reg [31:0] shiftedStoreDataQPreg_15; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_706;
  reg  addrKnownPReg_0; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_707;
  reg  addrKnownPReg_1; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_708;
  reg  addrKnownPReg_2; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_709;
  reg  addrKnownPReg_3; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_710;
  reg  addrKnownPReg_4; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_711;
  reg  addrKnownPReg_5; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_712;
  reg  addrKnownPReg_6; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_713;
  reg  addrKnownPReg_7; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_714;
  reg  addrKnownPReg_8; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_715;
  reg  addrKnownPReg_9; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_716;
  reg  addrKnownPReg_10; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_717;
  reg  addrKnownPReg_11; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_718;
  reg  addrKnownPReg_12; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_719;
  reg  addrKnownPReg_13; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_720;
  reg  addrKnownPReg_14; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_721;
  reg  addrKnownPReg_15; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_722;
  reg  dataKnownPReg_0; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_723;
  reg  dataKnownPReg_1; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_724;
  reg  dataKnownPReg_2; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_725;
  reg  dataKnownPReg_3; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_726;
  reg  dataKnownPReg_4; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_727;
  reg  dataKnownPReg_5; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_728;
  reg  dataKnownPReg_6; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_729;
  reg  dataKnownPReg_7; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_730;
  reg  dataKnownPReg_8; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_731;
  reg  dataKnownPReg_9; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_732;
  reg  dataKnownPReg_10; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_733;
  reg  dataKnownPReg_11; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_734;
  reg  dataKnownPReg_12; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_735;
  reg  dataKnownPReg_13; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_736;
  reg  dataKnownPReg_14; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_737;
  reg  dataKnownPReg_15; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_738;
  wire [1:0] _T_88276; // @[LoadQueue.scala 191:60:@35143.4]
  wire [1:0] _T_88277; // @[LoadQueue.scala 191:60:@35144.4]
  wire [2:0] _T_88278; // @[LoadQueue.scala 191:60:@35145.4]
  wire [2:0] _T_88279; // @[LoadQueue.scala 191:60:@35146.4]
  wire [2:0] _T_88280; // @[LoadQueue.scala 191:60:@35147.4]
  wire [2:0] _T_88281; // @[LoadQueue.scala 191:60:@35148.4]
  wire [3:0] _T_88282; // @[LoadQueue.scala 191:60:@35149.4]
  wire [3:0] _T_88283; // @[LoadQueue.scala 191:60:@35150.4]
  wire [3:0] _T_88284; // @[LoadQueue.scala 191:60:@35151.4]
  wire [3:0] _T_88285; // @[LoadQueue.scala 191:60:@35152.4]
  wire [3:0] _T_88286; // @[LoadQueue.scala 191:60:@35153.4]
  wire [3:0] _T_88287; // @[LoadQueue.scala 191:60:@35154.4]
  wire [3:0] _T_88288; // @[LoadQueue.scala 191:60:@35155.4]
  wire [3:0] _T_88289; // @[LoadQueue.scala 191:60:@35156.4]
  wire  _T_88292; // @[LoadQueue.scala 192:43:@35158.4]
  wire  _T_88293; // @[LoadQueue.scala 192:43:@35159.4]
  wire  _T_88294; // @[LoadQueue.scala 192:43:@35160.4]
  wire  _T_88295; // @[LoadQueue.scala 192:43:@35161.4]
  wire  _T_88296; // @[LoadQueue.scala 192:43:@35162.4]
  wire  _T_88297; // @[LoadQueue.scala 192:43:@35163.4]
  wire  _T_88298; // @[LoadQueue.scala 192:43:@35164.4]
  wire  _T_88299; // @[LoadQueue.scala 192:43:@35165.4]
  wire  _T_88300; // @[LoadQueue.scala 192:43:@35166.4]
  wire  _T_88301; // @[LoadQueue.scala 192:43:@35167.4]
  wire  _T_88302; // @[LoadQueue.scala 192:43:@35168.4]
  wire  _T_88303; // @[LoadQueue.scala 192:43:@35169.4]
  wire  _T_88304; // @[LoadQueue.scala 192:43:@35170.4]
  wire  _T_88305; // @[LoadQueue.scala 192:43:@35171.4]
  wire  _T_88306; // @[LoadQueue.scala 192:43:@35172.4]
  wire  _GEN_864; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_865; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_866; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_867; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_868; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_869; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_870; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_871; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_872; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_873; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_874; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_875; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_876; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_877; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_878; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_879; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_881; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_882; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_883; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_884; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_885; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_886; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_887; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_888; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_889; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_890; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_891; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_892; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_893; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_894; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_895; // @[LoadQueue.scala 194:31:@35175.6]
  wire [31:0] _GEN_897; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_898; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_899; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_900; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_901; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_902; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_903; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_904; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_905; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_906; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_907; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_908; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_909; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_910; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_911; // @[LoadQueue.scala 195:31:@35176.6]
  wire  lastConflict_0_0; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_1; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_2; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_3; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_4; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_5; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_6; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_7; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_8; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_9; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_10; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_11; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_12; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_13; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_14; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_15; // @[LoadQueue.scala 192:53:@35173.4]
  wire  canBypass_0; // @[LoadQueue.scala 192:53:@35173.4]
  wire [31:0] bypassVal_0; // @[LoadQueue.scala 192:53:@35173.4]
  wire [1:0] _T_88412; // @[LoadQueue.scala 191:60:@35230.4]
  wire [1:0] _T_88413; // @[LoadQueue.scala 191:60:@35231.4]
  wire [2:0] _T_88414; // @[LoadQueue.scala 191:60:@35232.4]
  wire [2:0] _T_88415; // @[LoadQueue.scala 191:60:@35233.4]
  wire [2:0] _T_88416; // @[LoadQueue.scala 191:60:@35234.4]
  wire [2:0] _T_88417; // @[LoadQueue.scala 191:60:@35235.4]
  wire [3:0] _T_88418; // @[LoadQueue.scala 191:60:@35236.4]
  wire [3:0] _T_88419; // @[LoadQueue.scala 191:60:@35237.4]
  wire [3:0] _T_88420; // @[LoadQueue.scala 191:60:@35238.4]
  wire [3:0] _T_88421; // @[LoadQueue.scala 191:60:@35239.4]
  wire [3:0] _T_88422; // @[LoadQueue.scala 191:60:@35240.4]
  wire [3:0] _T_88423; // @[LoadQueue.scala 191:60:@35241.4]
  wire [3:0] _T_88424; // @[LoadQueue.scala 191:60:@35242.4]
  wire [3:0] _T_88425; // @[LoadQueue.scala 191:60:@35243.4]
  wire  _T_88428; // @[LoadQueue.scala 192:43:@35245.4]
  wire  _T_88429; // @[LoadQueue.scala 192:43:@35246.4]
  wire  _T_88430; // @[LoadQueue.scala 192:43:@35247.4]
  wire  _T_88431; // @[LoadQueue.scala 192:43:@35248.4]
  wire  _T_88432; // @[LoadQueue.scala 192:43:@35249.4]
  wire  _T_88433; // @[LoadQueue.scala 192:43:@35250.4]
  wire  _T_88434; // @[LoadQueue.scala 192:43:@35251.4]
  wire  _T_88435; // @[LoadQueue.scala 192:43:@35252.4]
  wire  _T_88436; // @[LoadQueue.scala 192:43:@35253.4]
  wire  _T_88437; // @[LoadQueue.scala 192:43:@35254.4]
  wire  _T_88438; // @[LoadQueue.scala 192:43:@35255.4]
  wire  _T_88439; // @[LoadQueue.scala 192:43:@35256.4]
  wire  _T_88440; // @[LoadQueue.scala 192:43:@35257.4]
  wire  _T_88441; // @[LoadQueue.scala 192:43:@35258.4]
  wire  _T_88442; // @[LoadQueue.scala 192:43:@35259.4]
  wire  _GEN_930; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_931; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_932; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_933; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_934; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_935; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_936; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_937; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_938; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_939; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_940; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_941; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_942; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_943; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_944; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_945; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_947; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_948; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_949; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_950; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_951; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_952; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_953; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_954; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_955; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_956; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_957; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_958; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_959; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_960; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_961; // @[LoadQueue.scala 194:31:@35262.6]
  wire [31:0] _GEN_963; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_964; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_965; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_966; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_967; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_968; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_969; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_970; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_971; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_972; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_973; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_974; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_975; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_976; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_977; // @[LoadQueue.scala 195:31:@35263.6]
  wire  lastConflict_1_0; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_1; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_2; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_3; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_4; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_5; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_6; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_7; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_8; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_9; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_10; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_11; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_12; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_13; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_14; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_15; // @[LoadQueue.scala 192:53:@35260.4]
  wire  canBypass_1; // @[LoadQueue.scala 192:53:@35260.4]
  wire [31:0] bypassVal_1; // @[LoadQueue.scala 192:53:@35260.4]
  wire [1:0] _T_88548; // @[LoadQueue.scala 191:60:@35317.4]
  wire [1:0] _T_88549; // @[LoadQueue.scala 191:60:@35318.4]
  wire [2:0] _T_88550; // @[LoadQueue.scala 191:60:@35319.4]
  wire [2:0] _T_88551; // @[LoadQueue.scala 191:60:@35320.4]
  wire [2:0] _T_88552; // @[LoadQueue.scala 191:60:@35321.4]
  wire [2:0] _T_88553; // @[LoadQueue.scala 191:60:@35322.4]
  wire [3:0] _T_88554; // @[LoadQueue.scala 191:60:@35323.4]
  wire [3:0] _T_88555; // @[LoadQueue.scala 191:60:@35324.4]
  wire [3:0] _T_88556; // @[LoadQueue.scala 191:60:@35325.4]
  wire [3:0] _T_88557; // @[LoadQueue.scala 191:60:@35326.4]
  wire [3:0] _T_88558; // @[LoadQueue.scala 191:60:@35327.4]
  wire [3:0] _T_88559; // @[LoadQueue.scala 191:60:@35328.4]
  wire [3:0] _T_88560; // @[LoadQueue.scala 191:60:@35329.4]
  wire [3:0] _T_88561; // @[LoadQueue.scala 191:60:@35330.4]
  wire  _T_88564; // @[LoadQueue.scala 192:43:@35332.4]
  wire  _T_88565; // @[LoadQueue.scala 192:43:@35333.4]
  wire  _T_88566; // @[LoadQueue.scala 192:43:@35334.4]
  wire  _T_88567; // @[LoadQueue.scala 192:43:@35335.4]
  wire  _T_88568; // @[LoadQueue.scala 192:43:@35336.4]
  wire  _T_88569; // @[LoadQueue.scala 192:43:@35337.4]
  wire  _T_88570; // @[LoadQueue.scala 192:43:@35338.4]
  wire  _T_88571; // @[LoadQueue.scala 192:43:@35339.4]
  wire  _T_88572; // @[LoadQueue.scala 192:43:@35340.4]
  wire  _T_88573; // @[LoadQueue.scala 192:43:@35341.4]
  wire  _T_88574; // @[LoadQueue.scala 192:43:@35342.4]
  wire  _T_88575; // @[LoadQueue.scala 192:43:@35343.4]
  wire  _T_88576; // @[LoadQueue.scala 192:43:@35344.4]
  wire  _T_88577; // @[LoadQueue.scala 192:43:@35345.4]
  wire  _T_88578; // @[LoadQueue.scala 192:43:@35346.4]
  wire  _GEN_996; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_997; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_998; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_999; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1000; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1001; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1002; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1003; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1004; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1005; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1006; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1007; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1008; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1009; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1010; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1011; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1013; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1014; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1015; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1016; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1017; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1018; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1019; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1020; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1021; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1022; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1023; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1024; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1025; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1026; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1027; // @[LoadQueue.scala 194:31:@35349.6]
  wire [31:0] _GEN_1029; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1030; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1031; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1032; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1033; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1034; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1035; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1036; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1037; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1038; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1039; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1040; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1041; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1042; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1043; // @[LoadQueue.scala 195:31:@35350.6]
  wire  lastConflict_2_0; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_1; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_2; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_3; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_4; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_5; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_6; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_7; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_8; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_9; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_10; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_11; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_12; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_13; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_14; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_15; // @[LoadQueue.scala 192:53:@35347.4]
  wire  canBypass_2; // @[LoadQueue.scala 192:53:@35347.4]
  wire [31:0] bypassVal_2; // @[LoadQueue.scala 192:53:@35347.4]
  wire [1:0] _T_88684; // @[LoadQueue.scala 191:60:@35404.4]
  wire [1:0] _T_88685; // @[LoadQueue.scala 191:60:@35405.4]
  wire [2:0] _T_88686; // @[LoadQueue.scala 191:60:@35406.4]
  wire [2:0] _T_88687; // @[LoadQueue.scala 191:60:@35407.4]
  wire [2:0] _T_88688; // @[LoadQueue.scala 191:60:@35408.4]
  wire [2:0] _T_88689; // @[LoadQueue.scala 191:60:@35409.4]
  wire [3:0] _T_88690; // @[LoadQueue.scala 191:60:@35410.4]
  wire [3:0] _T_88691; // @[LoadQueue.scala 191:60:@35411.4]
  wire [3:0] _T_88692; // @[LoadQueue.scala 191:60:@35412.4]
  wire [3:0] _T_88693; // @[LoadQueue.scala 191:60:@35413.4]
  wire [3:0] _T_88694; // @[LoadQueue.scala 191:60:@35414.4]
  wire [3:0] _T_88695; // @[LoadQueue.scala 191:60:@35415.4]
  wire [3:0] _T_88696; // @[LoadQueue.scala 191:60:@35416.4]
  wire [3:0] _T_88697; // @[LoadQueue.scala 191:60:@35417.4]
  wire  _T_88700; // @[LoadQueue.scala 192:43:@35419.4]
  wire  _T_88701; // @[LoadQueue.scala 192:43:@35420.4]
  wire  _T_88702; // @[LoadQueue.scala 192:43:@35421.4]
  wire  _T_88703; // @[LoadQueue.scala 192:43:@35422.4]
  wire  _T_88704; // @[LoadQueue.scala 192:43:@35423.4]
  wire  _T_88705; // @[LoadQueue.scala 192:43:@35424.4]
  wire  _T_88706; // @[LoadQueue.scala 192:43:@35425.4]
  wire  _T_88707; // @[LoadQueue.scala 192:43:@35426.4]
  wire  _T_88708; // @[LoadQueue.scala 192:43:@35427.4]
  wire  _T_88709; // @[LoadQueue.scala 192:43:@35428.4]
  wire  _T_88710; // @[LoadQueue.scala 192:43:@35429.4]
  wire  _T_88711; // @[LoadQueue.scala 192:43:@35430.4]
  wire  _T_88712; // @[LoadQueue.scala 192:43:@35431.4]
  wire  _T_88713; // @[LoadQueue.scala 192:43:@35432.4]
  wire  _T_88714; // @[LoadQueue.scala 192:43:@35433.4]
  wire  _GEN_1062; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1063; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1064; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1065; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1066; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1067; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1068; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1069; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1070; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1071; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1072; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1073; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1074; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1075; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1076; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1077; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1079; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1080; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1081; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1082; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1083; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1084; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1085; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1086; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1087; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1088; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1089; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1090; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1091; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1092; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1093; // @[LoadQueue.scala 194:31:@35436.6]
  wire [31:0] _GEN_1095; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1096; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1097; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1098; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1099; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1100; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1101; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1102; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1103; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1104; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1105; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1106; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1107; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1108; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1109; // @[LoadQueue.scala 195:31:@35437.6]
  wire  lastConflict_3_0; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_1; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_2; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_3; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_4; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_5; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_6; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_7; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_8; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_9; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_10; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_11; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_12; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_13; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_14; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_15; // @[LoadQueue.scala 192:53:@35434.4]
  wire  canBypass_3; // @[LoadQueue.scala 192:53:@35434.4]
  wire [31:0] bypassVal_3; // @[LoadQueue.scala 192:53:@35434.4]
  wire [1:0] _T_88820; // @[LoadQueue.scala 191:60:@35491.4]
  wire [1:0] _T_88821; // @[LoadQueue.scala 191:60:@35492.4]
  wire [2:0] _T_88822; // @[LoadQueue.scala 191:60:@35493.4]
  wire [2:0] _T_88823; // @[LoadQueue.scala 191:60:@35494.4]
  wire [2:0] _T_88824; // @[LoadQueue.scala 191:60:@35495.4]
  wire [2:0] _T_88825; // @[LoadQueue.scala 191:60:@35496.4]
  wire [3:0] _T_88826; // @[LoadQueue.scala 191:60:@35497.4]
  wire [3:0] _T_88827; // @[LoadQueue.scala 191:60:@35498.4]
  wire [3:0] _T_88828; // @[LoadQueue.scala 191:60:@35499.4]
  wire [3:0] _T_88829; // @[LoadQueue.scala 191:60:@35500.4]
  wire [3:0] _T_88830; // @[LoadQueue.scala 191:60:@35501.4]
  wire [3:0] _T_88831; // @[LoadQueue.scala 191:60:@35502.4]
  wire [3:0] _T_88832; // @[LoadQueue.scala 191:60:@35503.4]
  wire [3:0] _T_88833; // @[LoadQueue.scala 191:60:@35504.4]
  wire  _T_88836; // @[LoadQueue.scala 192:43:@35506.4]
  wire  _T_88837; // @[LoadQueue.scala 192:43:@35507.4]
  wire  _T_88838; // @[LoadQueue.scala 192:43:@35508.4]
  wire  _T_88839; // @[LoadQueue.scala 192:43:@35509.4]
  wire  _T_88840; // @[LoadQueue.scala 192:43:@35510.4]
  wire  _T_88841; // @[LoadQueue.scala 192:43:@35511.4]
  wire  _T_88842; // @[LoadQueue.scala 192:43:@35512.4]
  wire  _T_88843; // @[LoadQueue.scala 192:43:@35513.4]
  wire  _T_88844; // @[LoadQueue.scala 192:43:@35514.4]
  wire  _T_88845; // @[LoadQueue.scala 192:43:@35515.4]
  wire  _T_88846; // @[LoadQueue.scala 192:43:@35516.4]
  wire  _T_88847; // @[LoadQueue.scala 192:43:@35517.4]
  wire  _T_88848; // @[LoadQueue.scala 192:43:@35518.4]
  wire  _T_88849; // @[LoadQueue.scala 192:43:@35519.4]
  wire  _T_88850; // @[LoadQueue.scala 192:43:@35520.4]
  wire  _GEN_1128; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1129; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1130; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1131; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1132; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1133; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1134; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1135; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1136; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1137; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1138; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1139; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1140; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1141; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1142; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1143; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1145; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1146; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1147; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1148; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1149; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1150; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1151; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1152; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1153; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1154; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1155; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1156; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1157; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1158; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1159; // @[LoadQueue.scala 194:31:@35523.6]
  wire [31:0] _GEN_1161; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1162; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1163; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1164; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1165; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1166; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1167; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1168; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1169; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1170; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1171; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1172; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1173; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1174; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1175; // @[LoadQueue.scala 195:31:@35524.6]
  wire  lastConflict_4_0; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_1; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_2; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_3; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_4; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_5; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_6; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_7; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_8; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_9; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_10; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_11; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_12; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_13; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_14; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_15; // @[LoadQueue.scala 192:53:@35521.4]
  wire  canBypass_4; // @[LoadQueue.scala 192:53:@35521.4]
  wire [31:0] bypassVal_4; // @[LoadQueue.scala 192:53:@35521.4]
  wire [1:0] _T_88956; // @[LoadQueue.scala 191:60:@35578.4]
  wire [1:0] _T_88957; // @[LoadQueue.scala 191:60:@35579.4]
  wire [2:0] _T_88958; // @[LoadQueue.scala 191:60:@35580.4]
  wire [2:0] _T_88959; // @[LoadQueue.scala 191:60:@35581.4]
  wire [2:0] _T_88960; // @[LoadQueue.scala 191:60:@35582.4]
  wire [2:0] _T_88961; // @[LoadQueue.scala 191:60:@35583.4]
  wire [3:0] _T_88962; // @[LoadQueue.scala 191:60:@35584.4]
  wire [3:0] _T_88963; // @[LoadQueue.scala 191:60:@35585.4]
  wire [3:0] _T_88964; // @[LoadQueue.scala 191:60:@35586.4]
  wire [3:0] _T_88965; // @[LoadQueue.scala 191:60:@35587.4]
  wire [3:0] _T_88966; // @[LoadQueue.scala 191:60:@35588.4]
  wire [3:0] _T_88967; // @[LoadQueue.scala 191:60:@35589.4]
  wire [3:0] _T_88968; // @[LoadQueue.scala 191:60:@35590.4]
  wire [3:0] _T_88969; // @[LoadQueue.scala 191:60:@35591.4]
  wire  _T_88972; // @[LoadQueue.scala 192:43:@35593.4]
  wire  _T_88973; // @[LoadQueue.scala 192:43:@35594.4]
  wire  _T_88974; // @[LoadQueue.scala 192:43:@35595.4]
  wire  _T_88975; // @[LoadQueue.scala 192:43:@35596.4]
  wire  _T_88976; // @[LoadQueue.scala 192:43:@35597.4]
  wire  _T_88977; // @[LoadQueue.scala 192:43:@35598.4]
  wire  _T_88978; // @[LoadQueue.scala 192:43:@35599.4]
  wire  _T_88979; // @[LoadQueue.scala 192:43:@35600.4]
  wire  _T_88980; // @[LoadQueue.scala 192:43:@35601.4]
  wire  _T_88981; // @[LoadQueue.scala 192:43:@35602.4]
  wire  _T_88982; // @[LoadQueue.scala 192:43:@35603.4]
  wire  _T_88983; // @[LoadQueue.scala 192:43:@35604.4]
  wire  _T_88984; // @[LoadQueue.scala 192:43:@35605.4]
  wire  _T_88985; // @[LoadQueue.scala 192:43:@35606.4]
  wire  _T_88986; // @[LoadQueue.scala 192:43:@35607.4]
  wire  _GEN_1194; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1195; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1196; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1197; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1198; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1199; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1200; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1201; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1202; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1203; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1204; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1205; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1206; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1207; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1208; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1209; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1211; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1212; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1213; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1214; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1215; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1216; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1217; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1218; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1219; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1220; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1221; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1222; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1223; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1224; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1225; // @[LoadQueue.scala 194:31:@35610.6]
  wire [31:0] _GEN_1227; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1228; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1229; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1230; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1231; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1232; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1233; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1234; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1235; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1236; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1237; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1238; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1239; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1240; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1241; // @[LoadQueue.scala 195:31:@35611.6]
  wire  lastConflict_5_0; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_1; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_2; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_3; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_4; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_5; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_6; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_7; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_8; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_9; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_10; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_11; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_12; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_13; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_14; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_15; // @[LoadQueue.scala 192:53:@35608.4]
  wire  canBypass_5; // @[LoadQueue.scala 192:53:@35608.4]
  wire [31:0] bypassVal_5; // @[LoadQueue.scala 192:53:@35608.4]
  wire [1:0] _T_89092; // @[LoadQueue.scala 191:60:@35665.4]
  wire [1:0] _T_89093; // @[LoadQueue.scala 191:60:@35666.4]
  wire [2:0] _T_89094; // @[LoadQueue.scala 191:60:@35667.4]
  wire [2:0] _T_89095; // @[LoadQueue.scala 191:60:@35668.4]
  wire [2:0] _T_89096; // @[LoadQueue.scala 191:60:@35669.4]
  wire [2:0] _T_89097; // @[LoadQueue.scala 191:60:@35670.4]
  wire [3:0] _T_89098; // @[LoadQueue.scala 191:60:@35671.4]
  wire [3:0] _T_89099; // @[LoadQueue.scala 191:60:@35672.4]
  wire [3:0] _T_89100; // @[LoadQueue.scala 191:60:@35673.4]
  wire [3:0] _T_89101; // @[LoadQueue.scala 191:60:@35674.4]
  wire [3:0] _T_89102; // @[LoadQueue.scala 191:60:@35675.4]
  wire [3:0] _T_89103; // @[LoadQueue.scala 191:60:@35676.4]
  wire [3:0] _T_89104; // @[LoadQueue.scala 191:60:@35677.4]
  wire [3:0] _T_89105; // @[LoadQueue.scala 191:60:@35678.4]
  wire  _T_89108; // @[LoadQueue.scala 192:43:@35680.4]
  wire  _T_89109; // @[LoadQueue.scala 192:43:@35681.4]
  wire  _T_89110; // @[LoadQueue.scala 192:43:@35682.4]
  wire  _T_89111; // @[LoadQueue.scala 192:43:@35683.4]
  wire  _T_89112; // @[LoadQueue.scala 192:43:@35684.4]
  wire  _T_89113; // @[LoadQueue.scala 192:43:@35685.4]
  wire  _T_89114; // @[LoadQueue.scala 192:43:@35686.4]
  wire  _T_89115; // @[LoadQueue.scala 192:43:@35687.4]
  wire  _T_89116; // @[LoadQueue.scala 192:43:@35688.4]
  wire  _T_89117; // @[LoadQueue.scala 192:43:@35689.4]
  wire  _T_89118; // @[LoadQueue.scala 192:43:@35690.4]
  wire  _T_89119; // @[LoadQueue.scala 192:43:@35691.4]
  wire  _T_89120; // @[LoadQueue.scala 192:43:@35692.4]
  wire  _T_89121; // @[LoadQueue.scala 192:43:@35693.4]
  wire  _T_89122; // @[LoadQueue.scala 192:43:@35694.4]
  wire  _GEN_1260; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1261; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1262; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1263; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1264; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1265; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1266; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1267; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1268; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1269; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1270; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1271; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1272; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1273; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1274; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1275; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1277; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1278; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1279; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1280; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1281; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1282; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1283; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1284; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1285; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1286; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1287; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1288; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1289; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1290; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1291; // @[LoadQueue.scala 194:31:@35697.6]
  wire [31:0] _GEN_1293; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1294; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1295; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1296; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1297; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1298; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1299; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1300; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1301; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1302; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1303; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1304; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1305; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1306; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1307; // @[LoadQueue.scala 195:31:@35698.6]
  wire  lastConflict_6_0; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_1; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_2; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_3; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_4; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_5; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_6; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_7; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_8; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_9; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_10; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_11; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_12; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_13; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_14; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_15; // @[LoadQueue.scala 192:53:@35695.4]
  wire  canBypass_6; // @[LoadQueue.scala 192:53:@35695.4]
  wire [31:0] bypassVal_6; // @[LoadQueue.scala 192:53:@35695.4]
  wire [1:0] _T_89228; // @[LoadQueue.scala 191:60:@35752.4]
  wire [1:0] _T_89229; // @[LoadQueue.scala 191:60:@35753.4]
  wire [2:0] _T_89230; // @[LoadQueue.scala 191:60:@35754.4]
  wire [2:0] _T_89231; // @[LoadQueue.scala 191:60:@35755.4]
  wire [2:0] _T_89232; // @[LoadQueue.scala 191:60:@35756.4]
  wire [2:0] _T_89233; // @[LoadQueue.scala 191:60:@35757.4]
  wire [3:0] _T_89234; // @[LoadQueue.scala 191:60:@35758.4]
  wire [3:0] _T_89235; // @[LoadQueue.scala 191:60:@35759.4]
  wire [3:0] _T_89236; // @[LoadQueue.scala 191:60:@35760.4]
  wire [3:0] _T_89237; // @[LoadQueue.scala 191:60:@35761.4]
  wire [3:0] _T_89238; // @[LoadQueue.scala 191:60:@35762.4]
  wire [3:0] _T_89239; // @[LoadQueue.scala 191:60:@35763.4]
  wire [3:0] _T_89240; // @[LoadQueue.scala 191:60:@35764.4]
  wire [3:0] _T_89241; // @[LoadQueue.scala 191:60:@35765.4]
  wire  _T_89244; // @[LoadQueue.scala 192:43:@35767.4]
  wire  _T_89245; // @[LoadQueue.scala 192:43:@35768.4]
  wire  _T_89246; // @[LoadQueue.scala 192:43:@35769.4]
  wire  _T_89247; // @[LoadQueue.scala 192:43:@35770.4]
  wire  _T_89248; // @[LoadQueue.scala 192:43:@35771.4]
  wire  _T_89249; // @[LoadQueue.scala 192:43:@35772.4]
  wire  _T_89250; // @[LoadQueue.scala 192:43:@35773.4]
  wire  _T_89251; // @[LoadQueue.scala 192:43:@35774.4]
  wire  _T_89252; // @[LoadQueue.scala 192:43:@35775.4]
  wire  _T_89253; // @[LoadQueue.scala 192:43:@35776.4]
  wire  _T_89254; // @[LoadQueue.scala 192:43:@35777.4]
  wire  _T_89255; // @[LoadQueue.scala 192:43:@35778.4]
  wire  _T_89256; // @[LoadQueue.scala 192:43:@35779.4]
  wire  _T_89257; // @[LoadQueue.scala 192:43:@35780.4]
  wire  _T_89258; // @[LoadQueue.scala 192:43:@35781.4]
  wire  _GEN_1326; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1327; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1328; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1329; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1330; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1331; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1332; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1333; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1334; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1335; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1336; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1337; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1338; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1339; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1340; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1341; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1343; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1344; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1345; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1346; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1347; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1348; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1349; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1350; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1351; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1352; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1353; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1354; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1355; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1356; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1357; // @[LoadQueue.scala 194:31:@35784.6]
  wire [31:0] _GEN_1359; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1360; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1361; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1362; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1363; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1364; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1365; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1366; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1367; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1368; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1369; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1370; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1371; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1372; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1373; // @[LoadQueue.scala 195:31:@35785.6]
  wire  lastConflict_7_0; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_1; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_2; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_3; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_4; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_5; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_6; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_7; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_8; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_9; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_10; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_11; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_12; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_13; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_14; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_15; // @[LoadQueue.scala 192:53:@35782.4]
  wire  canBypass_7; // @[LoadQueue.scala 192:53:@35782.4]
  wire [31:0] bypassVal_7; // @[LoadQueue.scala 192:53:@35782.4]
  wire [1:0] _T_89364; // @[LoadQueue.scala 191:60:@35839.4]
  wire [1:0] _T_89365; // @[LoadQueue.scala 191:60:@35840.4]
  wire [2:0] _T_89366; // @[LoadQueue.scala 191:60:@35841.4]
  wire [2:0] _T_89367; // @[LoadQueue.scala 191:60:@35842.4]
  wire [2:0] _T_89368; // @[LoadQueue.scala 191:60:@35843.4]
  wire [2:0] _T_89369; // @[LoadQueue.scala 191:60:@35844.4]
  wire [3:0] _T_89370; // @[LoadQueue.scala 191:60:@35845.4]
  wire [3:0] _T_89371; // @[LoadQueue.scala 191:60:@35846.4]
  wire [3:0] _T_89372; // @[LoadQueue.scala 191:60:@35847.4]
  wire [3:0] _T_89373; // @[LoadQueue.scala 191:60:@35848.4]
  wire [3:0] _T_89374; // @[LoadQueue.scala 191:60:@35849.4]
  wire [3:0] _T_89375; // @[LoadQueue.scala 191:60:@35850.4]
  wire [3:0] _T_89376; // @[LoadQueue.scala 191:60:@35851.4]
  wire [3:0] _T_89377; // @[LoadQueue.scala 191:60:@35852.4]
  wire  _T_89380; // @[LoadQueue.scala 192:43:@35854.4]
  wire  _T_89381; // @[LoadQueue.scala 192:43:@35855.4]
  wire  _T_89382; // @[LoadQueue.scala 192:43:@35856.4]
  wire  _T_89383; // @[LoadQueue.scala 192:43:@35857.4]
  wire  _T_89384; // @[LoadQueue.scala 192:43:@35858.4]
  wire  _T_89385; // @[LoadQueue.scala 192:43:@35859.4]
  wire  _T_89386; // @[LoadQueue.scala 192:43:@35860.4]
  wire  _T_89387; // @[LoadQueue.scala 192:43:@35861.4]
  wire  _T_89388; // @[LoadQueue.scala 192:43:@35862.4]
  wire  _T_89389; // @[LoadQueue.scala 192:43:@35863.4]
  wire  _T_89390; // @[LoadQueue.scala 192:43:@35864.4]
  wire  _T_89391; // @[LoadQueue.scala 192:43:@35865.4]
  wire  _T_89392; // @[LoadQueue.scala 192:43:@35866.4]
  wire  _T_89393; // @[LoadQueue.scala 192:43:@35867.4]
  wire  _T_89394; // @[LoadQueue.scala 192:43:@35868.4]
  wire  _GEN_1392; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1393; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1394; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1395; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1396; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1397; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1398; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1399; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1400; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1401; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1402; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1403; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1404; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1405; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1406; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1407; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1409; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1410; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1411; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1412; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1413; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1414; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1415; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1416; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1417; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1418; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1419; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1420; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1421; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1422; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1423; // @[LoadQueue.scala 194:31:@35871.6]
  wire [31:0] _GEN_1425; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1426; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1427; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1428; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1429; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1430; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1431; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1432; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1433; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1434; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1435; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1436; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1437; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1438; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1439; // @[LoadQueue.scala 195:31:@35872.6]
  wire  lastConflict_8_0; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_1; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_2; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_3; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_4; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_5; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_6; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_7; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_8; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_9; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_10; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_11; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_12; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_13; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_14; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_15; // @[LoadQueue.scala 192:53:@35869.4]
  wire  canBypass_8; // @[LoadQueue.scala 192:53:@35869.4]
  wire [31:0] bypassVal_8; // @[LoadQueue.scala 192:53:@35869.4]
  wire [1:0] _T_89500; // @[LoadQueue.scala 191:60:@35926.4]
  wire [1:0] _T_89501; // @[LoadQueue.scala 191:60:@35927.4]
  wire [2:0] _T_89502; // @[LoadQueue.scala 191:60:@35928.4]
  wire [2:0] _T_89503; // @[LoadQueue.scala 191:60:@35929.4]
  wire [2:0] _T_89504; // @[LoadQueue.scala 191:60:@35930.4]
  wire [2:0] _T_89505; // @[LoadQueue.scala 191:60:@35931.4]
  wire [3:0] _T_89506; // @[LoadQueue.scala 191:60:@35932.4]
  wire [3:0] _T_89507; // @[LoadQueue.scala 191:60:@35933.4]
  wire [3:0] _T_89508; // @[LoadQueue.scala 191:60:@35934.4]
  wire [3:0] _T_89509; // @[LoadQueue.scala 191:60:@35935.4]
  wire [3:0] _T_89510; // @[LoadQueue.scala 191:60:@35936.4]
  wire [3:0] _T_89511; // @[LoadQueue.scala 191:60:@35937.4]
  wire [3:0] _T_89512; // @[LoadQueue.scala 191:60:@35938.4]
  wire [3:0] _T_89513; // @[LoadQueue.scala 191:60:@35939.4]
  wire  _T_89516; // @[LoadQueue.scala 192:43:@35941.4]
  wire  _T_89517; // @[LoadQueue.scala 192:43:@35942.4]
  wire  _T_89518; // @[LoadQueue.scala 192:43:@35943.4]
  wire  _T_89519; // @[LoadQueue.scala 192:43:@35944.4]
  wire  _T_89520; // @[LoadQueue.scala 192:43:@35945.4]
  wire  _T_89521; // @[LoadQueue.scala 192:43:@35946.4]
  wire  _T_89522; // @[LoadQueue.scala 192:43:@35947.4]
  wire  _T_89523; // @[LoadQueue.scala 192:43:@35948.4]
  wire  _T_89524; // @[LoadQueue.scala 192:43:@35949.4]
  wire  _T_89525; // @[LoadQueue.scala 192:43:@35950.4]
  wire  _T_89526; // @[LoadQueue.scala 192:43:@35951.4]
  wire  _T_89527; // @[LoadQueue.scala 192:43:@35952.4]
  wire  _T_89528; // @[LoadQueue.scala 192:43:@35953.4]
  wire  _T_89529; // @[LoadQueue.scala 192:43:@35954.4]
  wire  _T_89530; // @[LoadQueue.scala 192:43:@35955.4]
  wire  _GEN_1458; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1459; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1460; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1461; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1462; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1463; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1464; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1465; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1466; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1467; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1468; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1469; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1470; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1471; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1472; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1473; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1475; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1476; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1477; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1478; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1479; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1480; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1481; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1482; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1483; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1484; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1485; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1486; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1487; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1488; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1489; // @[LoadQueue.scala 194:31:@35958.6]
  wire [31:0] _GEN_1491; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1492; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1493; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1494; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1495; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1496; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1497; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1498; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1499; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1500; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1501; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1502; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1503; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1504; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1505; // @[LoadQueue.scala 195:31:@35959.6]
  wire  lastConflict_9_0; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_1; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_2; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_3; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_4; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_5; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_6; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_7; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_8; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_9; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_10; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_11; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_12; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_13; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_14; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_15; // @[LoadQueue.scala 192:53:@35956.4]
  wire  canBypass_9; // @[LoadQueue.scala 192:53:@35956.4]
  wire [31:0] bypassVal_9; // @[LoadQueue.scala 192:53:@35956.4]
  wire [1:0] _T_89636; // @[LoadQueue.scala 191:60:@36013.4]
  wire [1:0] _T_89637; // @[LoadQueue.scala 191:60:@36014.4]
  wire [2:0] _T_89638; // @[LoadQueue.scala 191:60:@36015.4]
  wire [2:0] _T_89639; // @[LoadQueue.scala 191:60:@36016.4]
  wire [2:0] _T_89640; // @[LoadQueue.scala 191:60:@36017.4]
  wire [2:0] _T_89641; // @[LoadQueue.scala 191:60:@36018.4]
  wire [3:0] _T_89642; // @[LoadQueue.scala 191:60:@36019.4]
  wire [3:0] _T_89643; // @[LoadQueue.scala 191:60:@36020.4]
  wire [3:0] _T_89644; // @[LoadQueue.scala 191:60:@36021.4]
  wire [3:0] _T_89645; // @[LoadQueue.scala 191:60:@36022.4]
  wire [3:0] _T_89646; // @[LoadQueue.scala 191:60:@36023.4]
  wire [3:0] _T_89647; // @[LoadQueue.scala 191:60:@36024.4]
  wire [3:0] _T_89648; // @[LoadQueue.scala 191:60:@36025.4]
  wire [3:0] _T_89649; // @[LoadQueue.scala 191:60:@36026.4]
  wire  _T_89652; // @[LoadQueue.scala 192:43:@36028.4]
  wire  _T_89653; // @[LoadQueue.scala 192:43:@36029.4]
  wire  _T_89654; // @[LoadQueue.scala 192:43:@36030.4]
  wire  _T_89655; // @[LoadQueue.scala 192:43:@36031.4]
  wire  _T_89656; // @[LoadQueue.scala 192:43:@36032.4]
  wire  _T_89657; // @[LoadQueue.scala 192:43:@36033.4]
  wire  _T_89658; // @[LoadQueue.scala 192:43:@36034.4]
  wire  _T_89659; // @[LoadQueue.scala 192:43:@36035.4]
  wire  _T_89660; // @[LoadQueue.scala 192:43:@36036.4]
  wire  _T_89661; // @[LoadQueue.scala 192:43:@36037.4]
  wire  _T_89662; // @[LoadQueue.scala 192:43:@36038.4]
  wire  _T_89663; // @[LoadQueue.scala 192:43:@36039.4]
  wire  _T_89664; // @[LoadQueue.scala 192:43:@36040.4]
  wire  _T_89665; // @[LoadQueue.scala 192:43:@36041.4]
  wire  _T_89666; // @[LoadQueue.scala 192:43:@36042.4]
  wire  _GEN_1524; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1525; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1526; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1527; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1528; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1529; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1530; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1531; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1532; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1533; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1534; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1535; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1536; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1537; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1538; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1539; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1541; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1542; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1543; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1544; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1545; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1546; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1547; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1548; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1549; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1550; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1551; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1552; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1553; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1554; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1555; // @[LoadQueue.scala 194:31:@36045.6]
  wire [31:0] _GEN_1557; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1558; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1559; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1560; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1561; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1562; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1563; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1564; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1565; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1566; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1567; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1568; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1569; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1570; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1571; // @[LoadQueue.scala 195:31:@36046.6]
  wire  lastConflict_10_0; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_1; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_2; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_3; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_4; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_5; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_6; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_7; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_8; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_9; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_10; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_11; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_12; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_13; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_14; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_15; // @[LoadQueue.scala 192:53:@36043.4]
  wire  canBypass_10; // @[LoadQueue.scala 192:53:@36043.4]
  wire [31:0] bypassVal_10; // @[LoadQueue.scala 192:53:@36043.4]
  wire [1:0] _T_89772; // @[LoadQueue.scala 191:60:@36100.4]
  wire [1:0] _T_89773; // @[LoadQueue.scala 191:60:@36101.4]
  wire [2:0] _T_89774; // @[LoadQueue.scala 191:60:@36102.4]
  wire [2:0] _T_89775; // @[LoadQueue.scala 191:60:@36103.4]
  wire [2:0] _T_89776; // @[LoadQueue.scala 191:60:@36104.4]
  wire [2:0] _T_89777; // @[LoadQueue.scala 191:60:@36105.4]
  wire [3:0] _T_89778; // @[LoadQueue.scala 191:60:@36106.4]
  wire [3:0] _T_89779; // @[LoadQueue.scala 191:60:@36107.4]
  wire [3:0] _T_89780; // @[LoadQueue.scala 191:60:@36108.4]
  wire [3:0] _T_89781; // @[LoadQueue.scala 191:60:@36109.4]
  wire [3:0] _T_89782; // @[LoadQueue.scala 191:60:@36110.4]
  wire [3:0] _T_89783; // @[LoadQueue.scala 191:60:@36111.4]
  wire [3:0] _T_89784; // @[LoadQueue.scala 191:60:@36112.4]
  wire [3:0] _T_89785; // @[LoadQueue.scala 191:60:@36113.4]
  wire  _T_89788; // @[LoadQueue.scala 192:43:@36115.4]
  wire  _T_89789; // @[LoadQueue.scala 192:43:@36116.4]
  wire  _T_89790; // @[LoadQueue.scala 192:43:@36117.4]
  wire  _T_89791; // @[LoadQueue.scala 192:43:@36118.4]
  wire  _T_89792; // @[LoadQueue.scala 192:43:@36119.4]
  wire  _T_89793; // @[LoadQueue.scala 192:43:@36120.4]
  wire  _T_89794; // @[LoadQueue.scala 192:43:@36121.4]
  wire  _T_89795; // @[LoadQueue.scala 192:43:@36122.4]
  wire  _T_89796; // @[LoadQueue.scala 192:43:@36123.4]
  wire  _T_89797; // @[LoadQueue.scala 192:43:@36124.4]
  wire  _T_89798; // @[LoadQueue.scala 192:43:@36125.4]
  wire  _T_89799; // @[LoadQueue.scala 192:43:@36126.4]
  wire  _T_89800; // @[LoadQueue.scala 192:43:@36127.4]
  wire  _T_89801; // @[LoadQueue.scala 192:43:@36128.4]
  wire  _T_89802; // @[LoadQueue.scala 192:43:@36129.4]
  wire  _GEN_1590; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1591; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1592; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1593; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1594; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1595; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1596; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1597; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1598; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1599; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1600; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1601; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1602; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1603; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1604; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1605; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1607; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1608; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1609; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1610; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1611; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1612; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1613; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1614; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1615; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1616; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1617; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1618; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1619; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1620; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1621; // @[LoadQueue.scala 194:31:@36132.6]
  wire [31:0] _GEN_1623; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1624; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1625; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1626; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1627; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1628; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1629; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1630; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1631; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1632; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1633; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1634; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1635; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1636; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1637; // @[LoadQueue.scala 195:31:@36133.6]
  wire  lastConflict_11_0; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_1; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_2; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_3; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_4; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_5; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_6; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_7; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_8; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_9; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_10; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_11; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_12; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_13; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_14; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_15; // @[LoadQueue.scala 192:53:@36130.4]
  wire  canBypass_11; // @[LoadQueue.scala 192:53:@36130.4]
  wire [31:0] bypassVal_11; // @[LoadQueue.scala 192:53:@36130.4]
  wire [1:0] _T_89908; // @[LoadQueue.scala 191:60:@36187.4]
  wire [1:0] _T_89909; // @[LoadQueue.scala 191:60:@36188.4]
  wire [2:0] _T_89910; // @[LoadQueue.scala 191:60:@36189.4]
  wire [2:0] _T_89911; // @[LoadQueue.scala 191:60:@36190.4]
  wire [2:0] _T_89912; // @[LoadQueue.scala 191:60:@36191.4]
  wire [2:0] _T_89913; // @[LoadQueue.scala 191:60:@36192.4]
  wire [3:0] _T_89914; // @[LoadQueue.scala 191:60:@36193.4]
  wire [3:0] _T_89915; // @[LoadQueue.scala 191:60:@36194.4]
  wire [3:0] _T_89916; // @[LoadQueue.scala 191:60:@36195.4]
  wire [3:0] _T_89917; // @[LoadQueue.scala 191:60:@36196.4]
  wire [3:0] _T_89918; // @[LoadQueue.scala 191:60:@36197.4]
  wire [3:0] _T_89919; // @[LoadQueue.scala 191:60:@36198.4]
  wire [3:0] _T_89920; // @[LoadQueue.scala 191:60:@36199.4]
  wire [3:0] _T_89921; // @[LoadQueue.scala 191:60:@36200.4]
  wire  _T_89924; // @[LoadQueue.scala 192:43:@36202.4]
  wire  _T_89925; // @[LoadQueue.scala 192:43:@36203.4]
  wire  _T_89926; // @[LoadQueue.scala 192:43:@36204.4]
  wire  _T_89927; // @[LoadQueue.scala 192:43:@36205.4]
  wire  _T_89928; // @[LoadQueue.scala 192:43:@36206.4]
  wire  _T_89929; // @[LoadQueue.scala 192:43:@36207.4]
  wire  _T_89930; // @[LoadQueue.scala 192:43:@36208.4]
  wire  _T_89931; // @[LoadQueue.scala 192:43:@36209.4]
  wire  _T_89932; // @[LoadQueue.scala 192:43:@36210.4]
  wire  _T_89933; // @[LoadQueue.scala 192:43:@36211.4]
  wire  _T_89934; // @[LoadQueue.scala 192:43:@36212.4]
  wire  _T_89935; // @[LoadQueue.scala 192:43:@36213.4]
  wire  _T_89936; // @[LoadQueue.scala 192:43:@36214.4]
  wire  _T_89937; // @[LoadQueue.scala 192:43:@36215.4]
  wire  _T_89938; // @[LoadQueue.scala 192:43:@36216.4]
  wire  _GEN_1656; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1657; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1658; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1659; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1660; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1661; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1662; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1663; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1664; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1665; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1666; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1667; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1668; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1669; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1670; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1671; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1673; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1674; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1675; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1676; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1677; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1678; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1679; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1680; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1681; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1682; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1683; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1684; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1685; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1686; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1687; // @[LoadQueue.scala 194:31:@36219.6]
  wire [31:0] _GEN_1689; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1690; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1691; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1692; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1693; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1694; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1695; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1696; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1697; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1698; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1699; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1700; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1701; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1702; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1703; // @[LoadQueue.scala 195:31:@36220.6]
  wire  lastConflict_12_0; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_1; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_2; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_3; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_4; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_5; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_6; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_7; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_8; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_9; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_10; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_11; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_12; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_13; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_14; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_15; // @[LoadQueue.scala 192:53:@36217.4]
  wire  canBypass_12; // @[LoadQueue.scala 192:53:@36217.4]
  wire [31:0] bypassVal_12; // @[LoadQueue.scala 192:53:@36217.4]
  wire [1:0] _T_90044; // @[LoadQueue.scala 191:60:@36274.4]
  wire [1:0] _T_90045; // @[LoadQueue.scala 191:60:@36275.4]
  wire [2:0] _T_90046; // @[LoadQueue.scala 191:60:@36276.4]
  wire [2:0] _T_90047; // @[LoadQueue.scala 191:60:@36277.4]
  wire [2:0] _T_90048; // @[LoadQueue.scala 191:60:@36278.4]
  wire [2:0] _T_90049; // @[LoadQueue.scala 191:60:@36279.4]
  wire [3:0] _T_90050; // @[LoadQueue.scala 191:60:@36280.4]
  wire [3:0] _T_90051; // @[LoadQueue.scala 191:60:@36281.4]
  wire [3:0] _T_90052; // @[LoadQueue.scala 191:60:@36282.4]
  wire [3:0] _T_90053; // @[LoadQueue.scala 191:60:@36283.4]
  wire [3:0] _T_90054; // @[LoadQueue.scala 191:60:@36284.4]
  wire [3:0] _T_90055; // @[LoadQueue.scala 191:60:@36285.4]
  wire [3:0] _T_90056; // @[LoadQueue.scala 191:60:@36286.4]
  wire [3:0] _T_90057; // @[LoadQueue.scala 191:60:@36287.4]
  wire  _T_90060; // @[LoadQueue.scala 192:43:@36289.4]
  wire  _T_90061; // @[LoadQueue.scala 192:43:@36290.4]
  wire  _T_90062; // @[LoadQueue.scala 192:43:@36291.4]
  wire  _T_90063; // @[LoadQueue.scala 192:43:@36292.4]
  wire  _T_90064; // @[LoadQueue.scala 192:43:@36293.4]
  wire  _T_90065; // @[LoadQueue.scala 192:43:@36294.4]
  wire  _T_90066; // @[LoadQueue.scala 192:43:@36295.4]
  wire  _T_90067; // @[LoadQueue.scala 192:43:@36296.4]
  wire  _T_90068; // @[LoadQueue.scala 192:43:@36297.4]
  wire  _T_90069; // @[LoadQueue.scala 192:43:@36298.4]
  wire  _T_90070; // @[LoadQueue.scala 192:43:@36299.4]
  wire  _T_90071; // @[LoadQueue.scala 192:43:@36300.4]
  wire  _T_90072; // @[LoadQueue.scala 192:43:@36301.4]
  wire  _T_90073; // @[LoadQueue.scala 192:43:@36302.4]
  wire  _T_90074; // @[LoadQueue.scala 192:43:@36303.4]
  wire  _GEN_1722; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1723; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1724; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1725; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1726; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1727; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1728; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1729; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1730; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1731; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1732; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1733; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1734; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1735; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1736; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1737; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1739; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1740; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1741; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1742; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1743; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1744; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1745; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1746; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1747; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1748; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1749; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1750; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1751; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1752; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1753; // @[LoadQueue.scala 194:31:@36306.6]
  wire [31:0] _GEN_1755; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1756; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1757; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1758; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1759; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1760; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1761; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1762; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1763; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1764; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1765; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1766; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1767; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1768; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1769; // @[LoadQueue.scala 195:31:@36307.6]
  wire  lastConflict_13_0; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_1; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_2; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_3; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_4; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_5; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_6; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_7; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_8; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_9; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_10; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_11; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_12; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_13; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_14; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_15; // @[LoadQueue.scala 192:53:@36304.4]
  wire  canBypass_13; // @[LoadQueue.scala 192:53:@36304.4]
  wire [31:0] bypassVal_13; // @[LoadQueue.scala 192:53:@36304.4]
  wire [1:0] _T_90180; // @[LoadQueue.scala 191:60:@36361.4]
  wire [1:0] _T_90181; // @[LoadQueue.scala 191:60:@36362.4]
  wire [2:0] _T_90182; // @[LoadQueue.scala 191:60:@36363.4]
  wire [2:0] _T_90183; // @[LoadQueue.scala 191:60:@36364.4]
  wire [2:0] _T_90184; // @[LoadQueue.scala 191:60:@36365.4]
  wire [2:0] _T_90185; // @[LoadQueue.scala 191:60:@36366.4]
  wire [3:0] _T_90186; // @[LoadQueue.scala 191:60:@36367.4]
  wire [3:0] _T_90187; // @[LoadQueue.scala 191:60:@36368.4]
  wire [3:0] _T_90188; // @[LoadQueue.scala 191:60:@36369.4]
  wire [3:0] _T_90189; // @[LoadQueue.scala 191:60:@36370.4]
  wire [3:0] _T_90190; // @[LoadQueue.scala 191:60:@36371.4]
  wire [3:0] _T_90191; // @[LoadQueue.scala 191:60:@36372.4]
  wire [3:0] _T_90192; // @[LoadQueue.scala 191:60:@36373.4]
  wire [3:0] _T_90193; // @[LoadQueue.scala 191:60:@36374.4]
  wire  _T_90196; // @[LoadQueue.scala 192:43:@36376.4]
  wire  _T_90197; // @[LoadQueue.scala 192:43:@36377.4]
  wire  _T_90198; // @[LoadQueue.scala 192:43:@36378.4]
  wire  _T_90199; // @[LoadQueue.scala 192:43:@36379.4]
  wire  _T_90200; // @[LoadQueue.scala 192:43:@36380.4]
  wire  _T_90201; // @[LoadQueue.scala 192:43:@36381.4]
  wire  _T_90202; // @[LoadQueue.scala 192:43:@36382.4]
  wire  _T_90203; // @[LoadQueue.scala 192:43:@36383.4]
  wire  _T_90204; // @[LoadQueue.scala 192:43:@36384.4]
  wire  _T_90205; // @[LoadQueue.scala 192:43:@36385.4]
  wire  _T_90206; // @[LoadQueue.scala 192:43:@36386.4]
  wire  _T_90207; // @[LoadQueue.scala 192:43:@36387.4]
  wire  _T_90208; // @[LoadQueue.scala 192:43:@36388.4]
  wire  _T_90209; // @[LoadQueue.scala 192:43:@36389.4]
  wire  _T_90210; // @[LoadQueue.scala 192:43:@36390.4]
  wire  _GEN_1788; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1789; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1790; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1791; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1792; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1793; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1794; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1795; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1796; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1797; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1798; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1799; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1800; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1801; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1802; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1803; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1805; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1806; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1807; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1808; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1809; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1810; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1811; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1812; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1813; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1814; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1815; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1816; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1817; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1818; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1819; // @[LoadQueue.scala 194:31:@36393.6]
  wire [31:0] _GEN_1821; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1822; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1823; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1824; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1825; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1826; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1827; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1828; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1829; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1830; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1831; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1832; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1833; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1834; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1835; // @[LoadQueue.scala 195:31:@36394.6]
  wire  lastConflict_14_0; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_1; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_2; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_3; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_4; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_5; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_6; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_7; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_8; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_9; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_10; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_11; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_12; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_13; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_14; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_15; // @[LoadQueue.scala 192:53:@36391.4]
  wire  canBypass_14; // @[LoadQueue.scala 192:53:@36391.4]
  wire [31:0] bypassVal_14; // @[LoadQueue.scala 192:53:@36391.4]
  wire [1:0] _T_90316; // @[LoadQueue.scala 191:60:@36448.4]
  wire [1:0] _T_90317; // @[LoadQueue.scala 191:60:@36449.4]
  wire [2:0] _T_90318; // @[LoadQueue.scala 191:60:@36450.4]
  wire [2:0] _T_90319; // @[LoadQueue.scala 191:60:@36451.4]
  wire [2:0] _T_90320; // @[LoadQueue.scala 191:60:@36452.4]
  wire [2:0] _T_90321; // @[LoadQueue.scala 191:60:@36453.4]
  wire [3:0] _T_90322; // @[LoadQueue.scala 191:60:@36454.4]
  wire [3:0] _T_90323; // @[LoadQueue.scala 191:60:@36455.4]
  wire [3:0] _T_90324; // @[LoadQueue.scala 191:60:@36456.4]
  wire [3:0] _T_90325; // @[LoadQueue.scala 191:60:@36457.4]
  wire [3:0] _T_90326; // @[LoadQueue.scala 191:60:@36458.4]
  wire [3:0] _T_90327; // @[LoadQueue.scala 191:60:@36459.4]
  wire [3:0] _T_90328; // @[LoadQueue.scala 191:60:@36460.4]
  wire [3:0] _T_90329; // @[LoadQueue.scala 191:60:@36461.4]
  wire  _T_90332; // @[LoadQueue.scala 192:43:@36463.4]
  wire  _T_90333; // @[LoadQueue.scala 192:43:@36464.4]
  wire  _T_90334; // @[LoadQueue.scala 192:43:@36465.4]
  wire  _T_90335; // @[LoadQueue.scala 192:43:@36466.4]
  wire  _T_90336; // @[LoadQueue.scala 192:43:@36467.4]
  wire  _T_90337; // @[LoadQueue.scala 192:43:@36468.4]
  wire  _T_90338; // @[LoadQueue.scala 192:43:@36469.4]
  wire  _T_90339; // @[LoadQueue.scala 192:43:@36470.4]
  wire  _T_90340; // @[LoadQueue.scala 192:43:@36471.4]
  wire  _T_90341; // @[LoadQueue.scala 192:43:@36472.4]
  wire  _T_90342; // @[LoadQueue.scala 192:43:@36473.4]
  wire  _T_90343; // @[LoadQueue.scala 192:43:@36474.4]
  wire  _T_90344; // @[LoadQueue.scala 192:43:@36475.4]
  wire  _T_90345; // @[LoadQueue.scala 192:43:@36476.4]
  wire  _T_90346; // @[LoadQueue.scala 192:43:@36477.4]
  wire  _GEN_1854; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1855; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1856; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1857; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1858; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1859; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1860; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1861; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1862; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1863; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1864; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1865; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1866; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1867; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1868; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1869; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1871; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1872; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1873; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1874; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1875; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1876; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1877; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1878; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1879; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1880; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1881; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1882; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1883; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1884; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1885; // @[LoadQueue.scala 194:31:@36480.6]
  wire [31:0] _GEN_1887; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1888; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1889; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1890; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1891; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1892; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1893; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1894; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1895; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1896; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1897; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1898; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1899; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1900; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1901; // @[LoadQueue.scala 195:31:@36481.6]
  wire  lastConflict_15_0; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_1; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_2; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_3; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_4; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_5; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_6; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_7; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_8; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_9; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_10; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_11; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_12; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_13; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_14; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_15; // @[LoadQueue.scala 192:53:@36478.4]
  wire  canBypass_15; // @[LoadQueue.scala 192:53:@36478.4]
  wire [31:0] bypassVal_15; // @[LoadQueue.scala 192:53:@36478.4]
  wire [15:0] _T_90406; // @[OneHot.scala 52:12:@36486.4]
  wire  _T_90408; // @[util.scala 33:60:@36488.4]
  wire  _T_90409; // @[util.scala 33:60:@36489.4]
  wire  _T_90410; // @[util.scala 33:60:@36490.4]
  wire  _T_90411; // @[util.scala 33:60:@36491.4]
  wire  _T_90412; // @[util.scala 33:60:@36492.4]
  wire  _T_90413; // @[util.scala 33:60:@36493.4]
  wire  _T_90414; // @[util.scala 33:60:@36494.4]
  wire  _T_90415; // @[util.scala 33:60:@36495.4]
  wire  _T_90416; // @[util.scala 33:60:@36496.4]
  wire  _T_90417; // @[util.scala 33:60:@36497.4]
  wire  _T_90418; // @[util.scala 33:60:@36498.4]
  wire  _T_90419; // @[util.scala 33:60:@36499.4]
  wire  _T_90420; // @[util.scala 33:60:@36500.4]
  wire  _T_90421; // @[util.scala 33:60:@36501.4]
  wire  _T_90422; // @[util.scala 33:60:@36502.4]
  wire  _T_90423; // @[util.scala 33:60:@36503.4]
  wire  _T_93520; // @[LoadQueue.scala 229:41:@39026.4]
  wire  _T_93521; // @[LoadQueue.scala 229:38:@39027.4]
  wire  _T_93523; // @[LoadQueue.scala 230:12:@39029.6]
  reg  prevPriorityRequest_15; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_739;
  wire  _T_93525; // @[LoadQueue.scala 230:46:@39030.6]
  wire  _T_93526; // @[LoadQueue.scala 230:43:@39031.6]
  wire  _T_93528; // @[LoadQueue.scala 230:84:@39032.6]
  wire  _T_93529; // @[LoadQueue.scala 230:81:@39033.6]
  wire  _T_93532; // @[LoadQueue.scala 233:86:@39036.8]
  wire  _T_93533; // @[LoadQueue.scala 233:86:@39037.8]
  wire  _T_93534; // @[LoadQueue.scala 233:86:@39038.8]
  wire  _T_93535; // @[LoadQueue.scala 233:86:@39039.8]
  wire  _T_93536; // @[LoadQueue.scala 233:86:@39040.8]
  wire  _T_93537; // @[LoadQueue.scala 233:86:@39041.8]
  wire  _T_93538; // @[LoadQueue.scala 233:86:@39042.8]
  wire  _T_93539; // @[LoadQueue.scala 233:86:@39043.8]
  wire  _T_93540; // @[LoadQueue.scala 233:86:@39044.8]
  wire  _T_93541; // @[LoadQueue.scala 233:86:@39045.8]
  wire  _T_93542; // @[LoadQueue.scala 233:86:@39046.8]
  wire  _T_93543; // @[LoadQueue.scala 233:86:@39047.8]
  wire  _T_93544; // @[LoadQueue.scala 233:86:@39048.8]
  wire  _T_93545; // @[LoadQueue.scala 233:86:@39049.8]
  wire  _T_93546; // @[LoadQueue.scala 233:86:@39050.8]
  wire  _T_93548; // @[LoadQueue.scala 233:38:@39051.8]
  wire  _T_93567; // @[LoadQueue.scala 234:11:@39068.8]
  wire  _T_93568; // @[LoadQueue.scala 233:103:@39069.8]
  wire  _GEN_2028; // @[LoadQueue.scala 230:110:@39034.6]
  wire  loadRequest_15; // @[LoadQueue.scala 229:71:@39028.4]
  wire [15:0] _T_90464; // @[Mux.scala 31:69:@36521.4]
  wire  _T_93436; // @[LoadQueue.scala 229:41:@38944.4]
  wire  _T_93437; // @[LoadQueue.scala 229:38:@38945.4]
  wire  _T_93439; // @[LoadQueue.scala 230:12:@38947.6]
  reg  prevPriorityRequest_14; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_740;
  wire  _T_93441; // @[LoadQueue.scala 230:46:@38948.6]
  wire  _T_93442; // @[LoadQueue.scala 230:43:@38949.6]
  wire  _T_93444; // @[LoadQueue.scala 230:84:@38950.6]
  wire  _T_93445; // @[LoadQueue.scala 230:81:@38951.6]
  wire  _T_93448; // @[LoadQueue.scala 233:86:@38954.8]
  wire  _T_93449; // @[LoadQueue.scala 233:86:@38955.8]
  wire  _T_93450; // @[LoadQueue.scala 233:86:@38956.8]
  wire  _T_93451; // @[LoadQueue.scala 233:86:@38957.8]
  wire  _T_93452; // @[LoadQueue.scala 233:86:@38958.8]
  wire  _T_93453; // @[LoadQueue.scala 233:86:@38959.8]
  wire  _T_93454; // @[LoadQueue.scala 233:86:@38960.8]
  wire  _T_93455; // @[LoadQueue.scala 233:86:@38961.8]
  wire  _T_93456; // @[LoadQueue.scala 233:86:@38962.8]
  wire  _T_93457; // @[LoadQueue.scala 233:86:@38963.8]
  wire  _T_93458; // @[LoadQueue.scala 233:86:@38964.8]
  wire  _T_93459; // @[LoadQueue.scala 233:86:@38965.8]
  wire  _T_93460; // @[LoadQueue.scala 233:86:@38966.8]
  wire  _T_93461; // @[LoadQueue.scala 233:86:@38967.8]
  wire  _T_93462; // @[LoadQueue.scala 233:86:@38968.8]
  wire  _T_93464; // @[LoadQueue.scala 233:38:@38969.8]
  wire  _T_93483; // @[LoadQueue.scala 234:11:@38986.8]
  wire  _T_93484; // @[LoadQueue.scala 233:103:@38987.8]
  wire  _GEN_2024; // @[LoadQueue.scala 230:110:@38952.6]
  wire  loadRequest_14; // @[LoadQueue.scala 229:71:@38946.4]
  wire [15:0] _T_90465; // @[Mux.scala 31:69:@36522.4]
  wire  _T_93352; // @[LoadQueue.scala 229:41:@38862.4]
  wire  _T_93353; // @[LoadQueue.scala 229:38:@38863.4]
  wire  _T_93355; // @[LoadQueue.scala 230:12:@38865.6]
  reg  prevPriorityRequest_13; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_741;
  wire  _T_93357; // @[LoadQueue.scala 230:46:@38866.6]
  wire  _T_93358; // @[LoadQueue.scala 230:43:@38867.6]
  wire  _T_93360; // @[LoadQueue.scala 230:84:@38868.6]
  wire  _T_93361; // @[LoadQueue.scala 230:81:@38869.6]
  wire  _T_93364; // @[LoadQueue.scala 233:86:@38872.8]
  wire  _T_93365; // @[LoadQueue.scala 233:86:@38873.8]
  wire  _T_93366; // @[LoadQueue.scala 233:86:@38874.8]
  wire  _T_93367; // @[LoadQueue.scala 233:86:@38875.8]
  wire  _T_93368; // @[LoadQueue.scala 233:86:@38876.8]
  wire  _T_93369; // @[LoadQueue.scala 233:86:@38877.8]
  wire  _T_93370; // @[LoadQueue.scala 233:86:@38878.8]
  wire  _T_93371; // @[LoadQueue.scala 233:86:@38879.8]
  wire  _T_93372; // @[LoadQueue.scala 233:86:@38880.8]
  wire  _T_93373; // @[LoadQueue.scala 233:86:@38881.8]
  wire  _T_93374; // @[LoadQueue.scala 233:86:@38882.8]
  wire  _T_93375; // @[LoadQueue.scala 233:86:@38883.8]
  wire  _T_93376; // @[LoadQueue.scala 233:86:@38884.8]
  wire  _T_93377; // @[LoadQueue.scala 233:86:@38885.8]
  wire  _T_93378; // @[LoadQueue.scala 233:86:@38886.8]
  wire  _T_93380; // @[LoadQueue.scala 233:38:@38887.8]
  wire  _T_93399; // @[LoadQueue.scala 234:11:@38904.8]
  wire  _T_93400; // @[LoadQueue.scala 233:103:@38905.8]
  wire  _GEN_2020; // @[LoadQueue.scala 230:110:@38870.6]
  wire  loadRequest_13; // @[LoadQueue.scala 229:71:@38864.4]
  wire [15:0] _T_90466; // @[Mux.scala 31:69:@36523.4]
  wire  _T_93268; // @[LoadQueue.scala 229:41:@38780.4]
  wire  _T_93269; // @[LoadQueue.scala 229:38:@38781.4]
  wire  _T_93271; // @[LoadQueue.scala 230:12:@38783.6]
  reg  prevPriorityRequest_12; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_742;
  wire  _T_93273; // @[LoadQueue.scala 230:46:@38784.6]
  wire  _T_93274; // @[LoadQueue.scala 230:43:@38785.6]
  wire  _T_93276; // @[LoadQueue.scala 230:84:@38786.6]
  wire  _T_93277; // @[LoadQueue.scala 230:81:@38787.6]
  wire  _T_93280; // @[LoadQueue.scala 233:86:@38790.8]
  wire  _T_93281; // @[LoadQueue.scala 233:86:@38791.8]
  wire  _T_93282; // @[LoadQueue.scala 233:86:@38792.8]
  wire  _T_93283; // @[LoadQueue.scala 233:86:@38793.8]
  wire  _T_93284; // @[LoadQueue.scala 233:86:@38794.8]
  wire  _T_93285; // @[LoadQueue.scala 233:86:@38795.8]
  wire  _T_93286; // @[LoadQueue.scala 233:86:@38796.8]
  wire  _T_93287; // @[LoadQueue.scala 233:86:@38797.8]
  wire  _T_93288; // @[LoadQueue.scala 233:86:@38798.8]
  wire  _T_93289; // @[LoadQueue.scala 233:86:@38799.8]
  wire  _T_93290; // @[LoadQueue.scala 233:86:@38800.8]
  wire  _T_93291; // @[LoadQueue.scala 233:86:@38801.8]
  wire  _T_93292; // @[LoadQueue.scala 233:86:@38802.8]
  wire  _T_93293; // @[LoadQueue.scala 233:86:@38803.8]
  wire  _T_93294; // @[LoadQueue.scala 233:86:@38804.8]
  wire  _T_93296; // @[LoadQueue.scala 233:38:@38805.8]
  wire  _T_93315; // @[LoadQueue.scala 234:11:@38822.8]
  wire  _T_93316; // @[LoadQueue.scala 233:103:@38823.8]
  wire  _GEN_2016; // @[LoadQueue.scala 230:110:@38788.6]
  wire  loadRequest_12; // @[LoadQueue.scala 229:71:@38782.4]
  wire [15:0] _T_90467; // @[Mux.scala 31:69:@36524.4]
  wire  _T_93184; // @[LoadQueue.scala 229:41:@38698.4]
  wire  _T_93185; // @[LoadQueue.scala 229:38:@38699.4]
  wire  _T_93187; // @[LoadQueue.scala 230:12:@38701.6]
  reg  prevPriorityRequest_11; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_743;
  wire  _T_93189; // @[LoadQueue.scala 230:46:@38702.6]
  wire  _T_93190; // @[LoadQueue.scala 230:43:@38703.6]
  wire  _T_93192; // @[LoadQueue.scala 230:84:@38704.6]
  wire  _T_93193; // @[LoadQueue.scala 230:81:@38705.6]
  wire  _T_93196; // @[LoadQueue.scala 233:86:@38708.8]
  wire  _T_93197; // @[LoadQueue.scala 233:86:@38709.8]
  wire  _T_93198; // @[LoadQueue.scala 233:86:@38710.8]
  wire  _T_93199; // @[LoadQueue.scala 233:86:@38711.8]
  wire  _T_93200; // @[LoadQueue.scala 233:86:@38712.8]
  wire  _T_93201; // @[LoadQueue.scala 233:86:@38713.8]
  wire  _T_93202; // @[LoadQueue.scala 233:86:@38714.8]
  wire  _T_93203; // @[LoadQueue.scala 233:86:@38715.8]
  wire  _T_93204; // @[LoadQueue.scala 233:86:@38716.8]
  wire  _T_93205; // @[LoadQueue.scala 233:86:@38717.8]
  wire  _T_93206; // @[LoadQueue.scala 233:86:@38718.8]
  wire  _T_93207; // @[LoadQueue.scala 233:86:@38719.8]
  wire  _T_93208; // @[LoadQueue.scala 233:86:@38720.8]
  wire  _T_93209; // @[LoadQueue.scala 233:86:@38721.8]
  wire  _T_93210; // @[LoadQueue.scala 233:86:@38722.8]
  wire  _T_93212; // @[LoadQueue.scala 233:38:@38723.8]
  wire  _T_93231; // @[LoadQueue.scala 234:11:@38740.8]
  wire  _T_93232; // @[LoadQueue.scala 233:103:@38741.8]
  wire  _GEN_2012; // @[LoadQueue.scala 230:110:@38706.6]
  wire  loadRequest_11; // @[LoadQueue.scala 229:71:@38700.4]
  wire [15:0] _T_90468; // @[Mux.scala 31:69:@36525.4]
  wire  _T_93100; // @[LoadQueue.scala 229:41:@38616.4]
  wire  _T_93101; // @[LoadQueue.scala 229:38:@38617.4]
  wire  _T_93103; // @[LoadQueue.scala 230:12:@38619.6]
  reg  prevPriorityRequest_10; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_744;
  wire  _T_93105; // @[LoadQueue.scala 230:46:@38620.6]
  wire  _T_93106; // @[LoadQueue.scala 230:43:@38621.6]
  wire  _T_93108; // @[LoadQueue.scala 230:84:@38622.6]
  wire  _T_93109; // @[LoadQueue.scala 230:81:@38623.6]
  wire  _T_93112; // @[LoadQueue.scala 233:86:@38626.8]
  wire  _T_93113; // @[LoadQueue.scala 233:86:@38627.8]
  wire  _T_93114; // @[LoadQueue.scala 233:86:@38628.8]
  wire  _T_93115; // @[LoadQueue.scala 233:86:@38629.8]
  wire  _T_93116; // @[LoadQueue.scala 233:86:@38630.8]
  wire  _T_93117; // @[LoadQueue.scala 233:86:@38631.8]
  wire  _T_93118; // @[LoadQueue.scala 233:86:@38632.8]
  wire  _T_93119; // @[LoadQueue.scala 233:86:@38633.8]
  wire  _T_93120; // @[LoadQueue.scala 233:86:@38634.8]
  wire  _T_93121; // @[LoadQueue.scala 233:86:@38635.8]
  wire  _T_93122; // @[LoadQueue.scala 233:86:@38636.8]
  wire  _T_93123; // @[LoadQueue.scala 233:86:@38637.8]
  wire  _T_93124; // @[LoadQueue.scala 233:86:@38638.8]
  wire  _T_93125; // @[LoadQueue.scala 233:86:@38639.8]
  wire  _T_93126; // @[LoadQueue.scala 233:86:@38640.8]
  wire  _T_93128; // @[LoadQueue.scala 233:38:@38641.8]
  wire  _T_93147; // @[LoadQueue.scala 234:11:@38658.8]
  wire  _T_93148; // @[LoadQueue.scala 233:103:@38659.8]
  wire  _GEN_2008; // @[LoadQueue.scala 230:110:@38624.6]
  wire  loadRequest_10; // @[LoadQueue.scala 229:71:@38618.4]
  wire [15:0] _T_90469; // @[Mux.scala 31:69:@36526.4]
  wire  _T_93016; // @[LoadQueue.scala 229:41:@38534.4]
  wire  _T_93017; // @[LoadQueue.scala 229:38:@38535.4]
  wire  _T_93019; // @[LoadQueue.scala 230:12:@38537.6]
  reg  prevPriorityRequest_9; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_745;
  wire  _T_93021; // @[LoadQueue.scala 230:46:@38538.6]
  wire  _T_93022; // @[LoadQueue.scala 230:43:@38539.6]
  wire  _T_93024; // @[LoadQueue.scala 230:84:@38540.6]
  wire  _T_93025; // @[LoadQueue.scala 230:81:@38541.6]
  wire  _T_93028; // @[LoadQueue.scala 233:86:@38544.8]
  wire  _T_93029; // @[LoadQueue.scala 233:86:@38545.8]
  wire  _T_93030; // @[LoadQueue.scala 233:86:@38546.8]
  wire  _T_93031; // @[LoadQueue.scala 233:86:@38547.8]
  wire  _T_93032; // @[LoadQueue.scala 233:86:@38548.8]
  wire  _T_93033; // @[LoadQueue.scala 233:86:@38549.8]
  wire  _T_93034; // @[LoadQueue.scala 233:86:@38550.8]
  wire  _T_93035; // @[LoadQueue.scala 233:86:@38551.8]
  wire  _T_93036; // @[LoadQueue.scala 233:86:@38552.8]
  wire  _T_93037; // @[LoadQueue.scala 233:86:@38553.8]
  wire  _T_93038; // @[LoadQueue.scala 233:86:@38554.8]
  wire  _T_93039; // @[LoadQueue.scala 233:86:@38555.8]
  wire  _T_93040; // @[LoadQueue.scala 233:86:@38556.8]
  wire  _T_93041; // @[LoadQueue.scala 233:86:@38557.8]
  wire  _T_93042; // @[LoadQueue.scala 233:86:@38558.8]
  wire  _T_93044; // @[LoadQueue.scala 233:38:@38559.8]
  wire  _T_93063; // @[LoadQueue.scala 234:11:@38576.8]
  wire  _T_93064; // @[LoadQueue.scala 233:103:@38577.8]
  wire  _GEN_2004; // @[LoadQueue.scala 230:110:@38542.6]
  wire  loadRequest_9; // @[LoadQueue.scala 229:71:@38536.4]
  wire [15:0] _T_90470; // @[Mux.scala 31:69:@36527.4]
  wire  _T_92932; // @[LoadQueue.scala 229:41:@38452.4]
  wire  _T_92933; // @[LoadQueue.scala 229:38:@38453.4]
  wire  _T_92935; // @[LoadQueue.scala 230:12:@38455.6]
  reg  prevPriorityRequest_8; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_746;
  wire  _T_92937; // @[LoadQueue.scala 230:46:@38456.6]
  wire  _T_92938; // @[LoadQueue.scala 230:43:@38457.6]
  wire  _T_92940; // @[LoadQueue.scala 230:84:@38458.6]
  wire  _T_92941; // @[LoadQueue.scala 230:81:@38459.6]
  wire  _T_92944; // @[LoadQueue.scala 233:86:@38462.8]
  wire  _T_92945; // @[LoadQueue.scala 233:86:@38463.8]
  wire  _T_92946; // @[LoadQueue.scala 233:86:@38464.8]
  wire  _T_92947; // @[LoadQueue.scala 233:86:@38465.8]
  wire  _T_92948; // @[LoadQueue.scala 233:86:@38466.8]
  wire  _T_92949; // @[LoadQueue.scala 233:86:@38467.8]
  wire  _T_92950; // @[LoadQueue.scala 233:86:@38468.8]
  wire  _T_92951; // @[LoadQueue.scala 233:86:@38469.8]
  wire  _T_92952; // @[LoadQueue.scala 233:86:@38470.8]
  wire  _T_92953; // @[LoadQueue.scala 233:86:@38471.8]
  wire  _T_92954; // @[LoadQueue.scala 233:86:@38472.8]
  wire  _T_92955; // @[LoadQueue.scala 233:86:@38473.8]
  wire  _T_92956; // @[LoadQueue.scala 233:86:@38474.8]
  wire  _T_92957; // @[LoadQueue.scala 233:86:@38475.8]
  wire  _T_92958; // @[LoadQueue.scala 233:86:@38476.8]
  wire  _T_92960; // @[LoadQueue.scala 233:38:@38477.8]
  wire  _T_92979; // @[LoadQueue.scala 234:11:@38494.8]
  wire  _T_92980; // @[LoadQueue.scala 233:103:@38495.8]
  wire  _GEN_2000; // @[LoadQueue.scala 230:110:@38460.6]
  wire  loadRequest_8; // @[LoadQueue.scala 229:71:@38454.4]
  wire [15:0] _T_90471; // @[Mux.scala 31:69:@36528.4]
  wire  _T_92848; // @[LoadQueue.scala 229:41:@38370.4]
  wire  _T_92849; // @[LoadQueue.scala 229:38:@38371.4]
  wire  _T_92851; // @[LoadQueue.scala 230:12:@38373.6]
  reg  prevPriorityRequest_7; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_747;
  wire  _T_92853; // @[LoadQueue.scala 230:46:@38374.6]
  wire  _T_92854; // @[LoadQueue.scala 230:43:@38375.6]
  wire  _T_92856; // @[LoadQueue.scala 230:84:@38376.6]
  wire  _T_92857; // @[LoadQueue.scala 230:81:@38377.6]
  wire  _T_92860; // @[LoadQueue.scala 233:86:@38380.8]
  wire  _T_92861; // @[LoadQueue.scala 233:86:@38381.8]
  wire  _T_92862; // @[LoadQueue.scala 233:86:@38382.8]
  wire  _T_92863; // @[LoadQueue.scala 233:86:@38383.8]
  wire  _T_92864; // @[LoadQueue.scala 233:86:@38384.8]
  wire  _T_92865; // @[LoadQueue.scala 233:86:@38385.8]
  wire  _T_92866; // @[LoadQueue.scala 233:86:@38386.8]
  wire  _T_92867; // @[LoadQueue.scala 233:86:@38387.8]
  wire  _T_92868; // @[LoadQueue.scala 233:86:@38388.8]
  wire  _T_92869; // @[LoadQueue.scala 233:86:@38389.8]
  wire  _T_92870; // @[LoadQueue.scala 233:86:@38390.8]
  wire  _T_92871; // @[LoadQueue.scala 233:86:@38391.8]
  wire  _T_92872; // @[LoadQueue.scala 233:86:@38392.8]
  wire  _T_92873; // @[LoadQueue.scala 233:86:@38393.8]
  wire  _T_92874; // @[LoadQueue.scala 233:86:@38394.8]
  wire  _T_92876; // @[LoadQueue.scala 233:38:@38395.8]
  wire  _T_92895; // @[LoadQueue.scala 234:11:@38412.8]
  wire  _T_92896; // @[LoadQueue.scala 233:103:@38413.8]
  wire  _GEN_1996; // @[LoadQueue.scala 230:110:@38378.6]
  wire  loadRequest_7; // @[LoadQueue.scala 229:71:@38372.4]
  wire [15:0] _T_90472; // @[Mux.scala 31:69:@36529.4]
  wire  _T_92764; // @[LoadQueue.scala 229:41:@38288.4]
  wire  _T_92765; // @[LoadQueue.scala 229:38:@38289.4]
  wire  _T_92767; // @[LoadQueue.scala 230:12:@38291.6]
  reg  prevPriorityRequest_6; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_748;
  wire  _T_92769; // @[LoadQueue.scala 230:46:@38292.6]
  wire  _T_92770; // @[LoadQueue.scala 230:43:@38293.6]
  wire  _T_92772; // @[LoadQueue.scala 230:84:@38294.6]
  wire  _T_92773; // @[LoadQueue.scala 230:81:@38295.6]
  wire  _T_92776; // @[LoadQueue.scala 233:86:@38298.8]
  wire  _T_92777; // @[LoadQueue.scala 233:86:@38299.8]
  wire  _T_92778; // @[LoadQueue.scala 233:86:@38300.8]
  wire  _T_92779; // @[LoadQueue.scala 233:86:@38301.8]
  wire  _T_92780; // @[LoadQueue.scala 233:86:@38302.8]
  wire  _T_92781; // @[LoadQueue.scala 233:86:@38303.8]
  wire  _T_92782; // @[LoadQueue.scala 233:86:@38304.8]
  wire  _T_92783; // @[LoadQueue.scala 233:86:@38305.8]
  wire  _T_92784; // @[LoadQueue.scala 233:86:@38306.8]
  wire  _T_92785; // @[LoadQueue.scala 233:86:@38307.8]
  wire  _T_92786; // @[LoadQueue.scala 233:86:@38308.8]
  wire  _T_92787; // @[LoadQueue.scala 233:86:@38309.8]
  wire  _T_92788; // @[LoadQueue.scala 233:86:@38310.8]
  wire  _T_92789; // @[LoadQueue.scala 233:86:@38311.8]
  wire  _T_92790; // @[LoadQueue.scala 233:86:@38312.8]
  wire  _T_92792; // @[LoadQueue.scala 233:38:@38313.8]
  wire  _T_92811; // @[LoadQueue.scala 234:11:@38330.8]
  wire  _T_92812; // @[LoadQueue.scala 233:103:@38331.8]
  wire  _GEN_1992; // @[LoadQueue.scala 230:110:@38296.6]
  wire  loadRequest_6; // @[LoadQueue.scala 229:71:@38290.4]
  wire [15:0] _T_90473; // @[Mux.scala 31:69:@36530.4]
  wire  _T_92680; // @[LoadQueue.scala 229:41:@38206.4]
  wire  _T_92681; // @[LoadQueue.scala 229:38:@38207.4]
  wire  _T_92683; // @[LoadQueue.scala 230:12:@38209.6]
  reg  prevPriorityRequest_5; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_749;
  wire  _T_92685; // @[LoadQueue.scala 230:46:@38210.6]
  wire  _T_92686; // @[LoadQueue.scala 230:43:@38211.6]
  wire  _T_92688; // @[LoadQueue.scala 230:84:@38212.6]
  wire  _T_92689; // @[LoadQueue.scala 230:81:@38213.6]
  wire  _T_92692; // @[LoadQueue.scala 233:86:@38216.8]
  wire  _T_92693; // @[LoadQueue.scala 233:86:@38217.8]
  wire  _T_92694; // @[LoadQueue.scala 233:86:@38218.8]
  wire  _T_92695; // @[LoadQueue.scala 233:86:@38219.8]
  wire  _T_92696; // @[LoadQueue.scala 233:86:@38220.8]
  wire  _T_92697; // @[LoadQueue.scala 233:86:@38221.8]
  wire  _T_92698; // @[LoadQueue.scala 233:86:@38222.8]
  wire  _T_92699; // @[LoadQueue.scala 233:86:@38223.8]
  wire  _T_92700; // @[LoadQueue.scala 233:86:@38224.8]
  wire  _T_92701; // @[LoadQueue.scala 233:86:@38225.8]
  wire  _T_92702; // @[LoadQueue.scala 233:86:@38226.8]
  wire  _T_92703; // @[LoadQueue.scala 233:86:@38227.8]
  wire  _T_92704; // @[LoadQueue.scala 233:86:@38228.8]
  wire  _T_92705; // @[LoadQueue.scala 233:86:@38229.8]
  wire  _T_92706; // @[LoadQueue.scala 233:86:@38230.8]
  wire  _T_92708; // @[LoadQueue.scala 233:38:@38231.8]
  wire  _T_92727; // @[LoadQueue.scala 234:11:@38248.8]
  wire  _T_92728; // @[LoadQueue.scala 233:103:@38249.8]
  wire  _GEN_1988; // @[LoadQueue.scala 230:110:@38214.6]
  wire  loadRequest_5; // @[LoadQueue.scala 229:71:@38208.4]
  wire [15:0] _T_90474; // @[Mux.scala 31:69:@36531.4]
  wire  _T_92596; // @[LoadQueue.scala 229:41:@38124.4]
  wire  _T_92597; // @[LoadQueue.scala 229:38:@38125.4]
  wire  _T_92599; // @[LoadQueue.scala 230:12:@38127.6]
  reg  prevPriorityRequest_4; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_750;
  wire  _T_92601; // @[LoadQueue.scala 230:46:@38128.6]
  wire  _T_92602; // @[LoadQueue.scala 230:43:@38129.6]
  wire  _T_92604; // @[LoadQueue.scala 230:84:@38130.6]
  wire  _T_92605; // @[LoadQueue.scala 230:81:@38131.6]
  wire  _T_92608; // @[LoadQueue.scala 233:86:@38134.8]
  wire  _T_92609; // @[LoadQueue.scala 233:86:@38135.8]
  wire  _T_92610; // @[LoadQueue.scala 233:86:@38136.8]
  wire  _T_92611; // @[LoadQueue.scala 233:86:@38137.8]
  wire  _T_92612; // @[LoadQueue.scala 233:86:@38138.8]
  wire  _T_92613; // @[LoadQueue.scala 233:86:@38139.8]
  wire  _T_92614; // @[LoadQueue.scala 233:86:@38140.8]
  wire  _T_92615; // @[LoadQueue.scala 233:86:@38141.8]
  wire  _T_92616; // @[LoadQueue.scala 233:86:@38142.8]
  wire  _T_92617; // @[LoadQueue.scala 233:86:@38143.8]
  wire  _T_92618; // @[LoadQueue.scala 233:86:@38144.8]
  wire  _T_92619; // @[LoadQueue.scala 233:86:@38145.8]
  wire  _T_92620; // @[LoadQueue.scala 233:86:@38146.8]
  wire  _T_92621; // @[LoadQueue.scala 233:86:@38147.8]
  wire  _T_92622; // @[LoadQueue.scala 233:86:@38148.8]
  wire  _T_92624; // @[LoadQueue.scala 233:38:@38149.8]
  wire  _T_92643; // @[LoadQueue.scala 234:11:@38166.8]
  wire  _T_92644; // @[LoadQueue.scala 233:103:@38167.8]
  wire  _GEN_1984; // @[LoadQueue.scala 230:110:@38132.6]
  wire  loadRequest_4; // @[LoadQueue.scala 229:71:@38126.4]
  wire [15:0] _T_90475; // @[Mux.scala 31:69:@36532.4]
  wire  _T_92512; // @[LoadQueue.scala 229:41:@38042.4]
  wire  _T_92513; // @[LoadQueue.scala 229:38:@38043.4]
  wire  _T_92515; // @[LoadQueue.scala 230:12:@38045.6]
  reg  prevPriorityRequest_3; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_751;
  wire  _T_92517; // @[LoadQueue.scala 230:46:@38046.6]
  wire  _T_92518; // @[LoadQueue.scala 230:43:@38047.6]
  wire  _T_92520; // @[LoadQueue.scala 230:84:@38048.6]
  wire  _T_92521; // @[LoadQueue.scala 230:81:@38049.6]
  wire  _T_92524; // @[LoadQueue.scala 233:86:@38052.8]
  wire  _T_92525; // @[LoadQueue.scala 233:86:@38053.8]
  wire  _T_92526; // @[LoadQueue.scala 233:86:@38054.8]
  wire  _T_92527; // @[LoadQueue.scala 233:86:@38055.8]
  wire  _T_92528; // @[LoadQueue.scala 233:86:@38056.8]
  wire  _T_92529; // @[LoadQueue.scala 233:86:@38057.8]
  wire  _T_92530; // @[LoadQueue.scala 233:86:@38058.8]
  wire  _T_92531; // @[LoadQueue.scala 233:86:@38059.8]
  wire  _T_92532; // @[LoadQueue.scala 233:86:@38060.8]
  wire  _T_92533; // @[LoadQueue.scala 233:86:@38061.8]
  wire  _T_92534; // @[LoadQueue.scala 233:86:@38062.8]
  wire  _T_92535; // @[LoadQueue.scala 233:86:@38063.8]
  wire  _T_92536; // @[LoadQueue.scala 233:86:@38064.8]
  wire  _T_92537; // @[LoadQueue.scala 233:86:@38065.8]
  wire  _T_92538; // @[LoadQueue.scala 233:86:@38066.8]
  wire  _T_92540; // @[LoadQueue.scala 233:38:@38067.8]
  wire  _T_92559; // @[LoadQueue.scala 234:11:@38084.8]
  wire  _T_92560; // @[LoadQueue.scala 233:103:@38085.8]
  wire  _GEN_1980; // @[LoadQueue.scala 230:110:@38050.6]
  wire  loadRequest_3; // @[LoadQueue.scala 229:71:@38044.4]
  wire [15:0] _T_90476; // @[Mux.scala 31:69:@36533.4]
  wire  _T_92428; // @[LoadQueue.scala 229:41:@37960.4]
  wire  _T_92429; // @[LoadQueue.scala 229:38:@37961.4]
  wire  _T_92431; // @[LoadQueue.scala 230:12:@37963.6]
  reg  prevPriorityRequest_2; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_752;
  wire  _T_92433; // @[LoadQueue.scala 230:46:@37964.6]
  wire  _T_92434; // @[LoadQueue.scala 230:43:@37965.6]
  wire  _T_92436; // @[LoadQueue.scala 230:84:@37966.6]
  wire  _T_92437; // @[LoadQueue.scala 230:81:@37967.6]
  wire  _T_92440; // @[LoadQueue.scala 233:86:@37970.8]
  wire  _T_92441; // @[LoadQueue.scala 233:86:@37971.8]
  wire  _T_92442; // @[LoadQueue.scala 233:86:@37972.8]
  wire  _T_92443; // @[LoadQueue.scala 233:86:@37973.8]
  wire  _T_92444; // @[LoadQueue.scala 233:86:@37974.8]
  wire  _T_92445; // @[LoadQueue.scala 233:86:@37975.8]
  wire  _T_92446; // @[LoadQueue.scala 233:86:@37976.8]
  wire  _T_92447; // @[LoadQueue.scala 233:86:@37977.8]
  wire  _T_92448; // @[LoadQueue.scala 233:86:@37978.8]
  wire  _T_92449; // @[LoadQueue.scala 233:86:@37979.8]
  wire  _T_92450; // @[LoadQueue.scala 233:86:@37980.8]
  wire  _T_92451; // @[LoadQueue.scala 233:86:@37981.8]
  wire  _T_92452; // @[LoadQueue.scala 233:86:@37982.8]
  wire  _T_92453; // @[LoadQueue.scala 233:86:@37983.8]
  wire  _T_92454; // @[LoadQueue.scala 233:86:@37984.8]
  wire  _T_92456; // @[LoadQueue.scala 233:38:@37985.8]
  wire  _T_92475; // @[LoadQueue.scala 234:11:@38002.8]
  wire  _T_92476; // @[LoadQueue.scala 233:103:@38003.8]
  wire  _GEN_1976; // @[LoadQueue.scala 230:110:@37968.6]
  wire  loadRequest_2; // @[LoadQueue.scala 229:71:@37962.4]
  wire [15:0] _T_90477; // @[Mux.scala 31:69:@36534.4]
  wire  _T_92344; // @[LoadQueue.scala 229:41:@37878.4]
  wire  _T_92345; // @[LoadQueue.scala 229:38:@37879.4]
  wire  _T_92347; // @[LoadQueue.scala 230:12:@37881.6]
  reg  prevPriorityRequest_1; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_753;
  wire  _T_92349; // @[LoadQueue.scala 230:46:@37882.6]
  wire  _T_92350; // @[LoadQueue.scala 230:43:@37883.6]
  wire  _T_92352; // @[LoadQueue.scala 230:84:@37884.6]
  wire  _T_92353; // @[LoadQueue.scala 230:81:@37885.6]
  wire  _T_92356; // @[LoadQueue.scala 233:86:@37888.8]
  wire  _T_92357; // @[LoadQueue.scala 233:86:@37889.8]
  wire  _T_92358; // @[LoadQueue.scala 233:86:@37890.8]
  wire  _T_92359; // @[LoadQueue.scala 233:86:@37891.8]
  wire  _T_92360; // @[LoadQueue.scala 233:86:@37892.8]
  wire  _T_92361; // @[LoadQueue.scala 233:86:@37893.8]
  wire  _T_92362; // @[LoadQueue.scala 233:86:@37894.8]
  wire  _T_92363; // @[LoadQueue.scala 233:86:@37895.8]
  wire  _T_92364; // @[LoadQueue.scala 233:86:@37896.8]
  wire  _T_92365; // @[LoadQueue.scala 233:86:@37897.8]
  wire  _T_92366; // @[LoadQueue.scala 233:86:@37898.8]
  wire  _T_92367; // @[LoadQueue.scala 233:86:@37899.8]
  wire  _T_92368; // @[LoadQueue.scala 233:86:@37900.8]
  wire  _T_92369; // @[LoadQueue.scala 233:86:@37901.8]
  wire  _T_92370; // @[LoadQueue.scala 233:86:@37902.8]
  wire  _T_92372; // @[LoadQueue.scala 233:38:@37903.8]
  wire  _T_92391; // @[LoadQueue.scala 234:11:@37920.8]
  wire  _T_92392; // @[LoadQueue.scala 233:103:@37921.8]
  wire  _GEN_1972; // @[LoadQueue.scala 230:110:@37886.6]
  wire  loadRequest_1; // @[LoadQueue.scala 229:71:@37880.4]
  wire [15:0] _T_90478; // @[Mux.scala 31:69:@36535.4]
  wire  _T_92260; // @[LoadQueue.scala 229:41:@37796.4]
  wire  _T_92261; // @[LoadQueue.scala 229:38:@37797.4]
  wire  _T_92263; // @[LoadQueue.scala 230:12:@37799.6]
  reg  prevPriorityRequest_0; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_754;
  wire  _T_92265; // @[LoadQueue.scala 230:46:@37800.6]
  wire  _T_92266; // @[LoadQueue.scala 230:43:@37801.6]
  wire  _T_92268; // @[LoadQueue.scala 230:84:@37802.6]
  wire  _T_92269; // @[LoadQueue.scala 230:81:@37803.6]
  wire  _T_92272; // @[LoadQueue.scala 233:86:@37806.8]
  wire  _T_92273; // @[LoadQueue.scala 233:86:@37807.8]
  wire  _T_92274; // @[LoadQueue.scala 233:86:@37808.8]
  wire  _T_92275; // @[LoadQueue.scala 233:86:@37809.8]
  wire  _T_92276; // @[LoadQueue.scala 233:86:@37810.8]
  wire  _T_92277; // @[LoadQueue.scala 233:86:@37811.8]
  wire  _T_92278; // @[LoadQueue.scala 233:86:@37812.8]
  wire  _T_92279; // @[LoadQueue.scala 233:86:@37813.8]
  wire  _T_92280; // @[LoadQueue.scala 233:86:@37814.8]
  wire  _T_92281; // @[LoadQueue.scala 233:86:@37815.8]
  wire  _T_92282; // @[LoadQueue.scala 233:86:@37816.8]
  wire  _T_92283; // @[LoadQueue.scala 233:86:@37817.8]
  wire  _T_92284; // @[LoadQueue.scala 233:86:@37818.8]
  wire  _T_92285; // @[LoadQueue.scala 233:86:@37819.8]
  wire  _T_92286; // @[LoadQueue.scala 233:86:@37820.8]
  wire  _T_92288; // @[LoadQueue.scala 233:38:@37821.8]
  wire  _T_92307; // @[LoadQueue.scala 234:11:@37838.8]
  wire  _T_92308; // @[LoadQueue.scala 233:103:@37839.8]
  wire  _GEN_1968; // @[LoadQueue.scala 230:110:@37804.6]
  wire  loadRequest_0; // @[LoadQueue.scala 229:71:@37798.4]
  wire [15:0] _T_90479; // @[Mux.scala 31:69:@36536.4]
  wire  _T_90480; // @[OneHot.scala 66:30:@36537.4]
  wire  _T_90481; // @[OneHot.scala 66:30:@36538.4]
  wire  _T_90482; // @[OneHot.scala 66:30:@36539.4]
  wire  _T_90483; // @[OneHot.scala 66:30:@36540.4]
  wire  _T_90484; // @[OneHot.scala 66:30:@36541.4]
  wire  _T_90485; // @[OneHot.scala 66:30:@36542.4]
  wire  _T_90486; // @[OneHot.scala 66:30:@36543.4]
  wire  _T_90487; // @[OneHot.scala 66:30:@36544.4]
  wire  _T_90488; // @[OneHot.scala 66:30:@36545.4]
  wire  _T_90489; // @[OneHot.scala 66:30:@36546.4]
  wire  _T_90490; // @[OneHot.scala 66:30:@36547.4]
  wire  _T_90491; // @[OneHot.scala 66:30:@36548.4]
  wire  _T_90492; // @[OneHot.scala 66:30:@36549.4]
  wire  _T_90493; // @[OneHot.scala 66:30:@36550.4]
  wire  _T_90494; // @[OneHot.scala 66:30:@36551.4]
  wire  _T_90495; // @[OneHot.scala 66:30:@36552.4]
  wire [15:0] _T_90536; // @[Mux.scala 31:69:@36570.4]
  wire [15:0] _T_90537; // @[Mux.scala 31:69:@36571.4]
  wire [15:0] _T_90538; // @[Mux.scala 31:69:@36572.4]
  wire [15:0] _T_90539; // @[Mux.scala 31:69:@36573.4]
  wire [15:0] _T_90540; // @[Mux.scala 31:69:@36574.4]
  wire [15:0] _T_90541; // @[Mux.scala 31:69:@36575.4]
  wire [15:0] _T_90542; // @[Mux.scala 31:69:@36576.4]
  wire [15:0] _T_90543; // @[Mux.scala 31:69:@36577.4]
  wire [15:0] _T_90544; // @[Mux.scala 31:69:@36578.4]
  wire [15:0] _T_90545; // @[Mux.scala 31:69:@36579.4]
  wire [15:0] _T_90546; // @[Mux.scala 31:69:@36580.4]
  wire [15:0] _T_90547; // @[Mux.scala 31:69:@36581.4]
  wire [15:0] _T_90548; // @[Mux.scala 31:69:@36582.4]
  wire [15:0] _T_90549; // @[Mux.scala 31:69:@36583.4]
  wire [15:0] _T_90550; // @[Mux.scala 31:69:@36584.4]
  wire [15:0] _T_90551; // @[Mux.scala 31:69:@36585.4]
  wire  _T_90552; // @[OneHot.scala 66:30:@36586.4]
  wire  _T_90553; // @[OneHot.scala 66:30:@36587.4]
  wire  _T_90554; // @[OneHot.scala 66:30:@36588.4]
  wire  _T_90555; // @[OneHot.scala 66:30:@36589.4]
  wire  _T_90556; // @[OneHot.scala 66:30:@36590.4]
  wire  _T_90557; // @[OneHot.scala 66:30:@36591.4]
  wire  _T_90558; // @[OneHot.scala 66:30:@36592.4]
  wire  _T_90559; // @[OneHot.scala 66:30:@36593.4]
  wire  _T_90560; // @[OneHot.scala 66:30:@36594.4]
  wire  _T_90561; // @[OneHot.scala 66:30:@36595.4]
  wire  _T_90562; // @[OneHot.scala 66:30:@36596.4]
  wire  _T_90563; // @[OneHot.scala 66:30:@36597.4]
  wire  _T_90564; // @[OneHot.scala 66:30:@36598.4]
  wire  _T_90565; // @[OneHot.scala 66:30:@36599.4]
  wire  _T_90566; // @[OneHot.scala 66:30:@36600.4]
  wire  _T_90567; // @[OneHot.scala 66:30:@36601.4]
  wire [15:0] _T_90608; // @[Mux.scala 31:69:@36619.4]
  wire [15:0] _T_90609; // @[Mux.scala 31:69:@36620.4]
  wire [15:0] _T_90610; // @[Mux.scala 31:69:@36621.4]
  wire [15:0] _T_90611; // @[Mux.scala 31:69:@36622.4]
  wire [15:0] _T_90612; // @[Mux.scala 31:69:@36623.4]
  wire [15:0] _T_90613; // @[Mux.scala 31:69:@36624.4]
  wire [15:0] _T_90614; // @[Mux.scala 31:69:@36625.4]
  wire [15:0] _T_90615; // @[Mux.scala 31:69:@36626.4]
  wire [15:0] _T_90616; // @[Mux.scala 31:69:@36627.4]
  wire [15:0] _T_90617; // @[Mux.scala 31:69:@36628.4]
  wire [15:0] _T_90618; // @[Mux.scala 31:69:@36629.4]
  wire [15:0] _T_90619; // @[Mux.scala 31:69:@36630.4]
  wire [15:0] _T_90620; // @[Mux.scala 31:69:@36631.4]
  wire [15:0] _T_90621; // @[Mux.scala 31:69:@36632.4]
  wire [15:0] _T_90622; // @[Mux.scala 31:69:@36633.4]
  wire [15:0] _T_90623; // @[Mux.scala 31:69:@36634.4]
  wire  _T_90624; // @[OneHot.scala 66:30:@36635.4]
  wire  _T_90625; // @[OneHot.scala 66:30:@36636.4]
  wire  _T_90626; // @[OneHot.scala 66:30:@36637.4]
  wire  _T_90627; // @[OneHot.scala 66:30:@36638.4]
  wire  _T_90628; // @[OneHot.scala 66:30:@36639.4]
  wire  _T_90629; // @[OneHot.scala 66:30:@36640.4]
  wire  _T_90630; // @[OneHot.scala 66:30:@36641.4]
  wire  _T_90631; // @[OneHot.scala 66:30:@36642.4]
  wire  _T_90632; // @[OneHot.scala 66:30:@36643.4]
  wire  _T_90633; // @[OneHot.scala 66:30:@36644.4]
  wire  _T_90634; // @[OneHot.scala 66:30:@36645.4]
  wire  _T_90635; // @[OneHot.scala 66:30:@36646.4]
  wire  _T_90636; // @[OneHot.scala 66:30:@36647.4]
  wire  _T_90637; // @[OneHot.scala 66:30:@36648.4]
  wire  _T_90638; // @[OneHot.scala 66:30:@36649.4]
  wire  _T_90639; // @[OneHot.scala 66:30:@36650.4]
  wire [15:0] _T_90680; // @[Mux.scala 31:69:@36668.4]
  wire [15:0] _T_90681; // @[Mux.scala 31:69:@36669.4]
  wire [15:0] _T_90682; // @[Mux.scala 31:69:@36670.4]
  wire [15:0] _T_90683; // @[Mux.scala 31:69:@36671.4]
  wire [15:0] _T_90684; // @[Mux.scala 31:69:@36672.4]
  wire [15:0] _T_90685; // @[Mux.scala 31:69:@36673.4]
  wire [15:0] _T_90686; // @[Mux.scala 31:69:@36674.4]
  wire [15:0] _T_90687; // @[Mux.scala 31:69:@36675.4]
  wire [15:0] _T_90688; // @[Mux.scala 31:69:@36676.4]
  wire [15:0] _T_90689; // @[Mux.scala 31:69:@36677.4]
  wire [15:0] _T_90690; // @[Mux.scala 31:69:@36678.4]
  wire [15:0] _T_90691; // @[Mux.scala 31:69:@36679.4]
  wire [15:0] _T_90692; // @[Mux.scala 31:69:@36680.4]
  wire [15:0] _T_90693; // @[Mux.scala 31:69:@36681.4]
  wire [15:0] _T_90694; // @[Mux.scala 31:69:@36682.4]
  wire [15:0] _T_90695; // @[Mux.scala 31:69:@36683.4]
  wire  _T_90696; // @[OneHot.scala 66:30:@36684.4]
  wire  _T_90697; // @[OneHot.scala 66:30:@36685.4]
  wire  _T_90698; // @[OneHot.scala 66:30:@36686.4]
  wire  _T_90699; // @[OneHot.scala 66:30:@36687.4]
  wire  _T_90700; // @[OneHot.scala 66:30:@36688.4]
  wire  _T_90701; // @[OneHot.scala 66:30:@36689.4]
  wire  _T_90702; // @[OneHot.scala 66:30:@36690.4]
  wire  _T_90703; // @[OneHot.scala 66:30:@36691.4]
  wire  _T_90704; // @[OneHot.scala 66:30:@36692.4]
  wire  _T_90705; // @[OneHot.scala 66:30:@36693.4]
  wire  _T_90706; // @[OneHot.scala 66:30:@36694.4]
  wire  _T_90707; // @[OneHot.scala 66:30:@36695.4]
  wire  _T_90708; // @[OneHot.scala 66:30:@36696.4]
  wire  _T_90709; // @[OneHot.scala 66:30:@36697.4]
  wire  _T_90710; // @[OneHot.scala 66:30:@36698.4]
  wire  _T_90711; // @[OneHot.scala 66:30:@36699.4]
  wire [15:0] _T_90752; // @[Mux.scala 31:69:@36717.4]
  wire [15:0] _T_90753; // @[Mux.scala 31:69:@36718.4]
  wire [15:0] _T_90754; // @[Mux.scala 31:69:@36719.4]
  wire [15:0] _T_90755; // @[Mux.scala 31:69:@36720.4]
  wire [15:0] _T_90756; // @[Mux.scala 31:69:@36721.4]
  wire [15:0] _T_90757; // @[Mux.scala 31:69:@36722.4]
  wire [15:0] _T_90758; // @[Mux.scala 31:69:@36723.4]
  wire [15:0] _T_90759; // @[Mux.scala 31:69:@36724.4]
  wire [15:0] _T_90760; // @[Mux.scala 31:69:@36725.4]
  wire [15:0] _T_90761; // @[Mux.scala 31:69:@36726.4]
  wire [15:0] _T_90762; // @[Mux.scala 31:69:@36727.4]
  wire [15:0] _T_90763; // @[Mux.scala 31:69:@36728.4]
  wire [15:0] _T_90764; // @[Mux.scala 31:69:@36729.4]
  wire [15:0] _T_90765; // @[Mux.scala 31:69:@36730.4]
  wire [15:0] _T_90766; // @[Mux.scala 31:69:@36731.4]
  wire [15:0] _T_90767; // @[Mux.scala 31:69:@36732.4]
  wire  _T_90768; // @[OneHot.scala 66:30:@36733.4]
  wire  _T_90769; // @[OneHot.scala 66:30:@36734.4]
  wire  _T_90770; // @[OneHot.scala 66:30:@36735.4]
  wire  _T_90771; // @[OneHot.scala 66:30:@36736.4]
  wire  _T_90772; // @[OneHot.scala 66:30:@36737.4]
  wire  _T_90773; // @[OneHot.scala 66:30:@36738.4]
  wire  _T_90774; // @[OneHot.scala 66:30:@36739.4]
  wire  _T_90775; // @[OneHot.scala 66:30:@36740.4]
  wire  _T_90776; // @[OneHot.scala 66:30:@36741.4]
  wire  _T_90777; // @[OneHot.scala 66:30:@36742.4]
  wire  _T_90778; // @[OneHot.scala 66:30:@36743.4]
  wire  _T_90779; // @[OneHot.scala 66:30:@36744.4]
  wire  _T_90780; // @[OneHot.scala 66:30:@36745.4]
  wire  _T_90781; // @[OneHot.scala 66:30:@36746.4]
  wire  _T_90782; // @[OneHot.scala 66:30:@36747.4]
  wire  _T_90783; // @[OneHot.scala 66:30:@36748.4]
  wire [15:0] _T_90824; // @[Mux.scala 31:69:@36766.4]
  wire [15:0] _T_90825; // @[Mux.scala 31:69:@36767.4]
  wire [15:0] _T_90826; // @[Mux.scala 31:69:@36768.4]
  wire [15:0] _T_90827; // @[Mux.scala 31:69:@36769.4]
  wire [15:0] _T_90828; // @[Mux.scala 31:69:@36770.4]
  wire [15:0] _T_90829; // @[Mux.scala 31:69:@36771.4]
  wire [15:0] _T_90830; // @[Mux.scala 31:69:@36772.4]
  wire [15:0] _T_90831; // @[Mux.scala 31:69:@36773.4]
  wire [15:0] _T_90832; // @[Mux.scala 31:69:@36774.4]
  wire [15:0] _T_90833; // @[Mux.scala 31:69:@36775.4]
  wire [15:0] _T_90834; // @[Mux.scala 31:69:@36776.4]
  wire [15:0] _T_90835; // @[Mux.scala 31:69:@36777.4]
  wire [15:0] _T_90836; // @[Mux.scala 31:69:@36778.4]
  wire [15:0] _T_90837; // @[Mux.scala 31:69:@36779.4]
  wire [15:0] _T_90838; // @[Mux.scala 31:69:@36780.4]
  wire [15:0] _T_90839; // @[Mux.scala 31:69:@36781.4]
  wire  _T_90840; // @[OneHot.scala 66:30:@36782.4]
  wire  _T_90841; // @[OneHot.scala 66:30:@36783.4]
  wire  _T_90842; // @[OneHot.scala 66:30:@36784.4]
  wire  _T_90843; // @[OneHot.scala 66:30:@36785.4]
  wire  _T_90844; // @[OneHot.scala 66:30:@36786.4]
  wire  _T_90845; // @[OneHot.scala 66:30:@36787.4]
  wire  _T_90846; // @[OneHot.scala 66:30:@36788.4]
  wire  _T_90847; // @[OneHot.scala 66:30:@36789.4]
  wire  _T_90848; // @[OneHot.scala 66:30:@36790.4]
  wire  _T_90849; // @[OneHot.scala 66:30:@36791.4]
  wire  _T_90850; // @[OneHot.scala 66:30:@36792.4]
  wire  _T_90851; // @[OneHot.scala 66:30:@36793.4]
  wire  _T_90852; // @[OneHot.scala 66:30:@36794.4]
  wire  _T_90853; // @[OneHot.scala 66:30:@36795.4]
  wire  _T_90854; // @[OneHot.scala 66:30:@36796.4]
  wire  _T_90855; // @[OneHot.scala 66:30:@36797.4]
  wire [15:0] _T_90896; // @[Mux.scala 31:69:@36815.4]
  wire [15:0] _T_90897; // @[Mux.scala 31:69:@36816.4]
  wire [15:0] _T_90898; // @[Mux.scala 31:69:@36817.4]
  wire [15:0] _T_90899; // @[Mux.scala 31:69:@36818.4]
  wire [15:0] _T_90900; // @[Mux.scala 31:69:@36819.4]
  wire [15:0] _T_90901; // @[Mux.scala 31:69:@36820.4]
  wire [15:0] _T_90902; // @[Mux.scala 31:69:@36821.4]
  wire [15:0] _T_90903; // @[Mux.scala 31:69:@36822.4]
  wire [15:0] _T_90904; // @[Mux.scala 31:69:@36823.4]
  wire [15:0] _T_90905; // @[Mux.scala 31:69:@36824.4]
  wire [15:0] _T_90906; // @[Mux.scala 31:69:@36825.4]
  wire [15:0] _T_90907; // @[Mux.scala 31:69:@36826.4]
  wire [15:0] _T_90908; // @[Mux.scala 31:69:@36827.4]
  wire [15:0] _T_90909; // @[Mux.scala 31:69:@36828.4]
  wire [15:0] _T_90910; // @[Mux.scala 31:69:@36829.4]
  wire [15:0] _T_90911; // @[Mux.scala 31:69:@36830.4]
  wire  _T_90912; // @[OneHot.scala 66:30:@36831.4]
  wire  _T_90913; // @[OneHot.scala 66:30:@36832.4]
  wire  _T_90914; // @[OneHot.scala 66:30:@36833.4]
  wire  _T_90915; // @[OneHot.scala 66:30:@36834.4]
  wire  _T_90916; // @[OneHot.scala 66:30:@36835.4]
  wire  _T_90917; // @[OneHot.scala 66:30:@36836.4]
  wire  _T_90918; // @[OneHot.scala 66:30:@36837.4]
  wire  _T_90919; // @[OneHot.scala 66:30:@36838.4]
  wire  _T_90920; // @[OneHot.scala 66:30:@36839.4]
  wire  _T_90921; // @[OneHot.scala 66:30:@36840.4]
  wire  _T_90922; // @[OneHot.scala 66:30:@36841.4]
  wire  _T_90923; // @[OneHot.scala 66:30:@36842.4]
  wire  _T_90924; // @[OneHot.scala 66:30:@36843.4]
  wire  _T_90925; // @[OneHot.scala 66:30:@36844.4]
  wire  _T_90926; // @[OneHot.scala 66:30:@36845.4]
  wire  _T_90927; // @[OneHot.scala 66:30:@36846.4]
  wire [15:0] _T_90968; // @[Mux.scala 31:69:@36864.4]
  wire [15:0] _T_90969; // @[Mux.scala 31:69:@36865.4]
  wire [15:0] _T_90970; // @[Mux.scala 31:69:@36866.4]
  wire [15:0] _T_90971; // @[Mux.scala 31:69:@36867.4]
  wire [15:0] _T_90972; // @[Mux.scala 31:69:@36868.4]
  wire [15:0] _T_90973; // @[Mux.scala 31:69:@36869.4]
  wire [15:0] _T_90974; // @[Mux.scala 31:69:@36870.4]
  wire [15:0] _T_90975; // @[Mux.scala 31:69:@36871.4]
  wire [15:0] _T_90976; // @[Mux.scala 31:69:@36872.4]
  wire [15:0] _T_90977; // @[Mux.scala 31:69:@36873.4]
  wire [15:0] _T_90978; // @[Mux.scala 31:69:@36874.4]
  wire [15:0] _T_90979; // @[Mux.scala 31:69:@36875.4]
  wire [15:0] _T_90980; // @[Mux.scala 31:69:@36876.4]
  wire [15:0] _T_90981; // @[Mux.scala 31:69:@36877.4]
  wire [15:0] _T_90982; // @[Mux.scala 31:69:@36878.4]
  wire [15:0] _T_90983; // @[Mux.scala 31:69:@36879.4]
  wire  _T_90984; // @[OneHot.scala 66:30:@36880.4]
  wire  _T_90985; // @[OneHot.scala 66:30:@36881.4]
  wire  _T_90986; // @[OneHot.scala 66:30:@36882.4]
  wire  _T_90987; // @[OneHot.scala 66:30:@36883.4]
  wire  _T_90988; // @[OneHot.scala 66:30:@36884.4]
  wire  _T_90989; // @[OneHot.scala 66:30:@36885.4]
  wire  _T_90990; // @[OneHot.scala 66:30:@36886.4]
  wire  _T_90991; // @[OneHot.scala 66:30:@36887.4]
  wire  _T_90992; // @[OneHot.scala 66:30:@36888.4]
  wire  _T_90993; // @[OneHot.scala 66:30:@36889.4]
  wire  _T_90994; // @[OneHot.scala 66:30:@36890.4]
  wire  _T_90995; // @[OneHot.scala 66:30:@36891.4]
  wire  _T_90996; // @[OneHot.scala 66:30:@36892.4]
  wire  _T_90997; // @[OneHot.scala 66:30:@36893.4]
  wire  _T_90998; // @[OneHot.scala 66:30:@36894.4]
  wire  _T_90999; // @[OneHot.scala 66:30:@36895.4]
  wire [15:0] _T_91040; // @[Mux.scala 31:69:@36913.4]
  wire [15:0] _T_91041; // @[Mux.scala 31:69:@36914.4]
  wire [15:0] _T_91042; // @[Mux.scala 31:69:@36915.4]
  wire [15:0] _T_91043; // @[Mux.scala 31:69:@36916.4]
  wire [15:0] _T_91044; // @[Mux.scala 31:69:@36917.4]
  wire [15:0] _T_91045; // @[Mux.scala 31:69:@36918.4]
  wire [15:0] _T_91046; // @[Mux.scala 31:69:@36919.4]
  wire [15:0] _T_91047; // @[Mux.scala 31:69:@36920.4]
  wire [15:0] _T_91048; // @[Mux.scala 31:69:@36921.4]
  wire [15:0] _T_91049; // @[Mux.scala 31:69:@36922.4]
  wire [15:0] _T_91050; // @[Mux.scala 31:69:@36923.4]
  wire [15:0] _T_91051; // @[Mux.scala 31:69:@36924.4]
  wire [15:0] _T_91052; // @[Mux.scala 31:69:@36925.4]
  wire [15:0] _T_91053; // @[Mux.scala 31:69:@36926.4]
  wire [15:0] _T_91054; // @[Mux.scala 31:69:@36927.4]
  wire [15:0] _T_91055; // @[Mux.scala 31:69:@36928.4]
  wire  _T_91056; // @[OneHot.scala 66:30:@36929.4]
  wire  _T_91057; // @[OneHot.scala 66:30:@36930.4]
  wire  _T_91058; // @[OneHot.scala 66:30:@36931.4]
  wire  _T_91059; // @[OneHot.scala 66:30:@36932.4]
  wire  _T_91060; // @[OneHot.scala 66:30:@36933.4]
  wire  _T_91061; // @[OneHot.scala 66:30:@36934.4]
  wire  _T_91062; // @[OneHot.scala 66:30:@36935.4]
  wire  _T_91063; // @[OneHot.scala 66:30:@36936.4]
  wire  _T_91064; // @[OneHot.scala 66:30:@36937.4]
  wire  _T_91065; // @[OneHot.scala 66:30:@36938.4]
  wire  _T_91066; // @[OneHot.scala 66:30:@36939.4]
  wire  _T_91067; // @[OneHot.scala 66:30:@36940.4]
  wire  _T_91068; // @[OneHot.scala 66:30:@36941.4]
  wire  _T_91069; // @[OneHot.scala 66:30:@36942.4]
  wire  _T_91070; // @[OneHot.scala 66:30:@36943.4]
  wire  _T_91071; // @[OneHot.scala 66:30:@36944.4]
  wire [15:0] _T_91112; // @[Mux.scala 31:69:@36962.4]
  wire [15:0] _T_91113; // @[Mux.scala 31:69:@36963.4]
  wire [15:0] _T_91114; // @[Mux.scala 31:69:@36964.4]
  wire [15:0] _T_91115; // @[Mux.scala 31:69:@36965.4]
  wire [15:0] _T_91116; // @[Mux.scala 31:69:@36966.4]
  wire [15:0] _T_91117; // @[Mux.scala 31:69:@36967.4]
  wire [15:0] _T_91118; // @[Mux.scala 31:69:@36968.4]
  wire [15:0] _T_91119; // @[Mux.scala 31:69:@36969.4]
  wire [15:0] _T_91120; // @[Mux.scala 31:69:@36970.4]
  wire [15:0] _T_91121; // @[Mux.scala 31:69:@36971.4]
  wire [15:0] _T_91122; // @[Mux.scala 31:69:@36972.4]
  wire [15:0] _T_91123; // @[Mux.scala 31:69:@36973.4]
  wire [15:0] _T_91124; // @[Mux.scala 31:69:@36974.4]
  wire [15:0] _T_91125; // @[Mux.scala 31:69:@36975.4]
  wire [15:0] _T_91126; // @[Mux.scala 31:69:@36976.4]
  wire [15:0] _T_91127; // @[Mux.scala 31:69:@36977.4]
  wire  _T_91128; // @[OneHot.scala 66:30:@36978.4]
  wire  _T_91129; // @[OneHot.scala 66:30:@36979.4]
  wire  _T_91130; // @[OneHot.scala 66:30:@36980.4]
  wire  _T_91131; // @[OneHot.scala 66:30:@36981.4]
  wire  _T_91132; // @[OneHot.scala 66:30:@36982.4]
  wire  _T_91133; // @[OneHot.scala 66:30:@36983.4]
  wire  _T_91134; // @[OneHot.scala 66:30:@36984.4]
  wire  _T_91135; // @[OneHot.scala 66:30:@36985.4]
  wire  _T_91136; // @[OneHot.scala 66:30:@36986.4]
  wire  _T_91137; // @[OneHot.scala 66:30:@36987.4]
  wire  _T_91138; // @[OneHot.scala 66:30:@36988.4]
  wire  _T_91139; // @[OneHot.scala 66:30:@36989.4]
  wire  _T_91140; // @[OneHot.scala 66:30:@36990.4]
  wire  _T_91141; // @[OneHot.scala 66:30:@36991.4]
  wire  _T_91142; // @[OneHot.scala 66:30:@36992.4]
  wire  _T_91143; // @[OneHot.scala 66:30:@36993.4]
  wire [15:0] _T_91184; // @[Mux.scala 31:69:@37011.4]
  wire [15:0] _T_91185; // @[Mux.scala 31:69:@37012.4]
  wire [15:0] _T_91186; // @[Mux.scala 31:69:@37013.4]
  wire [15:0] _T_91187; // @[Mux.scala 31:69:@37014.4]
  wire [15:0] _T_91188; // @[Mux.scala 31:69:@37015.4]
  wire [15:0] _T_91189; // @[Mux.scala 31:69:@37016.4]
  wire [15:0] _T_91190; // @[Mux.scala 31:69:@37017.4]
  wire [15:0] _T_91191; // @[Mux.scala 31:69:@37018.4]
  wire [15:0] _T_91192; // @[Mux.scala 31:69:@37019.4]
  wire [15:0] _T_91193; // @[Mux.scala 31:69:@37020.4]
  wire [15:0] _T_91194; // @[Mux.scala 31:69:@37021.4]
  wire [15:0] _T_91195; // @[Mux.scala 31:69:@37022.4]
  wire [15:0] _T_91196; // @[Mux.scala 31:69:@37023.4]
  wire [15:0] _T_91197; // @[Mux.scala 31:69:@37024.4]
  wire [15:0] _T_91198; // @[Mux.scala 31:69:@37025.4]
  wire [15:0] _T_91199; // @[Mux.scala 31:69:@37026.4]
  wire  _T_91200; // @[OneHot.scala 66:30:@37027.4]
  wire  _T_91201; // @[OneHot.scala 66:30:@37028.4]
  wire  _T_91202; // @[OneHot.scala 66:30:@37029.4]
  wire  _T_91203; // @[OneHot.scala 66:30:@37030.4]
  wire  _T_91204; // @[OneHot.scala 66:30:@37031.4]
  wire  _T_91205; // @[OneHot.scala 66:30:@37032.4]
  wire  _T_91206; // @[OneHot.scala 66:30:@37033.4]
  wire  _T_91207; // @[OneHot.scala 66:30:@37034.4]
  wire  _T_91208; // @[OneHot.scala 66:30:@37035.4]
  wire  _T_91209; // @[OneHot.scala 66:30:@37036.4]
  wire  _T_91210; // @[OneHot.scala 66:30:@37037.4]
  wire  _T_91211; // @[OneHot.scala 66:30:@37038.4]
  wire  _T_91212; // @[OneHot.scala 66:30:@37039.4]
  wire  _T_91213; // @[OneHot.scala 66:30:@37040.4]
  wire  _T_91214; // @[OneHot.scala 66:30:@37041.4]
  wire  _T_91215; // @[OneHot.scala 66:30:@37042.4]
  wire [15:0] _T_91256; // @[Mux.scala 31:69:@37060.4]
  wire [15:0] _T_91257; // @[Mux.scala 31:69:@37061.4]
  wire [15:0] _T_91258; // @[Mux.scala 31:69:@37062.4]
  wire [15:0] _T_91259; // @[Mux.scala 31:69:@37063.4]
  wire [15:0] _T_91260; // @[Mux.scala 31:69:@37064.4]
  wire [15:0] _T_91261; // @[Mux.scala 31:69:@37065.4]
  wire [15:0] _T_91262; // @[Mux.scala 31:69:@37066.4]
  wire [15:0] _T_91263; // @[Mux.scala 31:69:@37067.4]
  wire [15:0] _T_91264; // @[Mux.scala 31:69:@37068.4]
  wire [15:0] _T_91265; // @[Mux.scala 31:69:@37069.4]
  wire [15:0] _T_91266; // @[Mux.scala 31:69:@37070.4]
  wire [15:0] _T_91267; // @[Mux.scala 31:69:@37071.4]
  wire [15:0] _T_91268; // @[Mux.scala 31:69:@37072.4]
  wire [15:0] _T_91269; // @[Mux.scala 31:69:@37073.4]
  wire [15:0] _T_91270; // @[Mux.scala 31:69:@37074.4]
  wire [15:0] _T_91271; // @[Mux.scala 31:69:@37075.4]
  wire  _T_91272; // @[OneHot.scala 66:30:@37076.4]
  wire  _T_91273; // @[OneHot.scala 66:30:@37077.4]
  wire  _T_91274; // @[OneHot.scala 66:30:@37078.4]
  wire  _T_91275; // @[OneHot.scala 66:30:@37079.4]
  wire  _T_91276; // @[OneHot.scala 66:30:@37080.4]
  wire  _T_91277; // @[OneHot.scala 66:30:@37081.4]
  wire  _T_91278; // @[OneHot.scala 66:30:@37082.4]
  wire  _T_91279; // @[OneHot.scala 66:30:@37083.4]
  wire  _T_91280; // @[OneHot.scala 66:30:@37084.4]
  wire  _T_91281; // @[OneHot.scala 66:30:@37085.4]
  wire  _T_91282; // @[OneHot.scala 66:30:@37086.4]
  wire  _T_91283; // @[OneHot.scala 66:30:@37087.4]
  wire  _T_91284; // @[OneHot.scala 66:30:@37088.4]
  wire  _T_91285; // @[OneHot.scala 66:30:@37089.4]
  wire  _T_91286; // @[OneHot.scala 66:30:@37090.4]
  wire  _T_91287; // @[OneHot.scala 66:30:@37091.4]
  wire [15:0] _T_91328; // @[Mux.scala 31:69:@37109.4]
  wire [15:0] _T_91329; // @[Mux.scala 31:69:@37110.4]
  wire [15:0] _T_91330; // @[Mux.scala 31:69:@37111.4]
  wire [15:0] _T_91331; // @[Mux.scala 31:69:@37112.4]
  wire [15:0] _T_91332; // @[Mux.scala 31:69:@37113.4]
  wire [15:0] _T_91333; // @[Mux.scala 31:69:@37114.4]
  wire [15:0] _T_91334; // @[Mux.scala 31:69:@37115.4]
  wire [15:0] _T_91335; // @[Mux.scala 31:69:@37116.4]
  wire [15:0] _T_91336; // @[Mux.scala 31:69:@37117.4]
  wire [15:0] _T_91337; // @[Mux.scala 31:69:@37118.4]
  wire [15:0] _T_91338; // @[Mux.scala 31:69:@37119.4]
  wire [15:0] _T_91339; // @[Mux.scala 31:69:@37120.4]
  wire [15:0] _T_91340; // @[Mux.scala 31:69:@37121.4]
  wire [15:0] _T_91341; // @[Mux.scala 31:69:@37122.4]
  wire [15:0] _T_91342; // @[Mux.scala 31:69:@37123.4]
  wire [15:0] _T_91343; // @[Mux.scala 31:69:@37124.4]
  wire  _T_91344; // @[OneHot.scala 66:30:@37125.4]
  wire  _T_91345; // @[OneHot.scala 66:30:@37126.4]
  wire  _T_91346; // @[OneHot.scala 66:30:@37127.4]
  wire  _T_91347; // @[OneHot.scala 66:30:@37128.4]
  wire  _T_91348; // @[OneHot.scala 66:30:@37129.4]
  wire  _T_91349; // @[OneHot.scala 66:30:@37130.4]
  wire  _T_91350; // @[OneHot.scala 66:30:@37131.4]
  wire  _T_91351; // @[OneHot.scala 66:30:@37132.4]
  wire  _T_91352; // @[OneHot.scala 66:30:@37133.4]
  wire  _T_91353; // @[OneHot.scala 66:30:@37134.4]
  wire  _T_91354; // @[OneHot.scala 66:30:@37135.4]
  wire  _T_91355; // @[OneHot.scala 66:30:@37136.4]
  wire  _T_91356; // @[OneHot.scala 66:30:@37137.4]
  wire  _T_91357; // @[OneHot.scala 66:30:@37138.4]
  wire  _T_91358; // @[OneHot.scala 66:30:@37139.4]
  wire  _T_91359; // @[OneHot.scala 66:30:@37140.4]
  wire [15:0] _T_91400; // @[Mux.scala 31:69:@37158.4]
  wire [15:0] _T_91401; // @[Mux.scala 31:69:@37159.4]
  wire [15:0] _T_91402; // @[Mux.scala 31:69:@37160.4]
  wire [15:0] _T_91403; // @[Mux.scala 31:69:@37161.4]
  wire [15:0] _T_91404; // @[Mux.scala 31:69:@37162.4]
  wire [15:0] _T_91405; // @[Mux.scala 31:69:@37163.4]
  wire [15:0] _T_91406; // @[Mux.scala 31:69:@37164.4]
  wire [15:0] _T_91407; // @[Mux.scala 31:69:@37165.4]
  wire [15:0] _T_91408; // @[Mux.scala 31:69:@37166.4]
  wire [15:0] _T_91409; // @[Mux.scala 31:69:@37167.4]
  wire [15:0] _T_91410; // @[Mux.scala 31:69:@37168.4]
  wire [15:0] _T_91411; // @[Mux.scala 31:69:@37169.4]
  wire [15:0] _T_91412; // @[Mux.scala 31:69:@37170.4]
  wire [15:0] _T_91413; // @[Mux.scala 31:69:@37171.4]
  wire [15:0] _T_91414; // @[Mux.scala 31:69:@37172.4]
  wire [15:0] _T_91415; // @[Mux.scala 31:69:@37173.4]
  wire  _T_91416; // @[OneHot.scala 66:30:@37174.4]
  wire  _T_91417; // @[OneHot.scala 66:30:@37175.4]
  wire  _T_91418; // @[OneHot.scala 66:30:@37176.4]
  wire  _T_91419; // @[OneHot.scala 66:30:@37177.4]
  wire  _T_91420; // @[OneHot.scala 66:30:@37178.4]
  wire  _T_91421; // @[OneHot.scala 66:30:@37179.4]
  wire  _T_91422; // @[OneHot.scala 66:30:@37180.4]
  wire  _T_91423; // @[OneHot.scala 66:30:@37181.4]
  wire  _T_91424; // @[OneHot.scala 66:30:@37182.4]
  wire  _T_91425; // @[OneHot.scala 66:30:@37183.4]
  wire  _T_91426; // @[OneHot.scala 66:30:@37184.4]
  wire  _T_91427; // @[OneHot.scala 66:30:@37185.4]
  wire  _T_91428; // @[OneHot.scala 66:30:@37186.4]
  wire  _T_91429; // @[OneHot.scala 66:30:@37187.4]
  wire  _T_91430; // @[OneHot.scala 66:30:@37188.4]
  wire  _T_91431; // @[OneHot.scala 66:30:@37189.4]
  wire [15:0] _T_91472; // @[Mux.scala 31:69:@37207.4]
  wire [15:0] _T_91473; // @[Mux.scala 31:69:@37208.4]
  wire [15:0] _T_91474; // @[Mux.scala 31:69:@37209.4]
  wire [15:0] _T_91475; // @[Mux.scala 31:69:@37210.4]
  wire [15:0] _T_91476; // @[Mux.scala 31:69:@37211.4]
  wire [15:0] _T_91477; // @[Mux.scala 31:69:@37212.4]
  wire [15:0] _T_91478; // @[Mux.scala 31:69:@37213.4]
  wire [15:0] _T_91479; // @[Mux.scala 31:69:@37214.4]
  wire [15:0] _T_91480; // @[Mux.scala 31:69:@37215.4]
  wire [15:0] _T_91481; // @[Mux.scala 31:69:@37216.4]
  wire [15:0] _T_91482; // @[Mux.scala 31:69:@37217.4]
  wire [15:0] _T_91483; // @[Mux.scala 31:69:@37218.4]
  wire [15:0] _T_91484; // @[Mux.scala 31:69:@37219.4]
  wire [15:0] _T_91485; // @[Mux.scala 31:69:@37220.4]
  wire [15:0] _T_91486; // @[Mux.scala 31:69:@37221.4]
  wire [15:0] _T_91487; // @[Mux.scala 31:69:@37222.4]
  wire  _T_91488; // @[OneHot.scala 66:30:@37223.4]
  wire  _T_91489; // @[OneHot.scala 66:30:@37224.4]
  wire  _T_91490; // @[OneHot.scala 66:30:@37225.4]
  wire  _T_91491; // @[OneHot.scala 66:30:@37226.4]
  wire  _T_91492; // @[OneHot.scala 66:30:@37227.4]
  wire  _T_91493; // @[OneHot.scala 66:30:@37228.4]
  wire  _T_91494; // @[OneHot.scala 66:30:@37229.4]
  wire  _T_91495; // @[OneHot.scala 66:30:@37230.4]
  wire  _T_91496; // @[OneHot.scala 66:30:@37231.4]
  wire  _T_91497; // @[OneHot.scala 66:30:@37232.4]
  wire  _T_91498; // @[OneHot.scala 66:30:@37233.4]
  wire  _T_91499; // @[OneHot.scala 66:30:@37234.4]
  wire  _T_91500; // @[OneHot.scala 66:30:@37235.4]
  wire  _T_91501; // @[OneHot.scala 66:30:@37236.4]
  wire  _T_91502; // @[OneHot.scala 66:30:@37237.4]
  wire  _T_91503; // @[OneHot.scala 66:30:@37238.4]
  wire [15:0] _T_91544; // @[Mux.scala 31:69:@37256.4]
  wire [15:0] _T_91545; // @[Mux.scala 31:69:@37257.4]
  wire [15:0] _T_91546; // @[Mux.scala 31:69:@37258.4]
  wire [15:0] _T_91547; // @[Mux.scala 31:69:@37259.4]
  wire [15:0] _T_91548; // @[Mux.scala 31:69:@37260.4]
  wire [15:0] _T_91549; // @[Mux.scala 31:69:@37261.4]
  wire [15:0] _T_91550; // @[Mux.scala 31:69:@37262.4]
  wire [15:0] _T_91551; // @[Mux.scala 31:69:@37263.4]
  wire [15:0] _T_91552; // @[Mux.scala 31:69:@37264.4]
  wire [15:0] _T_91553; // @[Mux.scala 31:69:@37265.4]
  wire [15:0] _T_91554; // @[Mux.scala 31:69:@37266.4]
  wire [15:0] _T_91555; // @[Mux.scala 31:69:@37267.4]
  wire [15:0] _T_91556; // @[Mux.scala 31:69:@37268.4]
  wire [15:0] _T_91557; // @[Mux.scala 31:69:@37269.4]
  wire [15:0] _T_91558; // @[Mux.scala 31:69:@37270.4]
  wire [15:0] _T_91559; // @[Mux.scala 31:69:@37271.4]
  wire  _T_91560; // @[OneHot.scala 66:30:@37272.4]
  wire  _T_91561; // @[OneHot.scala 66:30:@37273.4]
  wire  _T_91562; // @[OneHot.scala 66:30:@37274.4]
  wire  _T_91563; // @[OneHot.scala 66:30:@37275.4]
  wire  _T_91564; // @[OneHot.scala 66:30:@37276.4]
  wire  _T_91565; // @[OneHot.scala 66:30:@37277.4]
  wire  _T_91566; // @[OneHot.scala 66:30:@37278.4]
  wire  _T_91567; // @[OneHot.scala 66:30:@37279.4]
  wire  _T_91568; // @[OneHot.scala 66:30:@37280.4]
  wire  _T_91569; // @[OneHot.scala 66:30:@37281.4]
  wire  _T_91570; // @[OneHot.scala 66:30:@37282.4]
  wire  _T_91571; // @[OneHot.scala 66:30:@37283.4]
  wire  _T_91572; // @[OneHot.scala 66:30:@37284.4]
  wire  _T_91573; // @[OneHot.scala 66:30:@37285.4]
  wire  _T_91574; // @[OneHot.scala 66:30:@37286.4]
  wire  _T_91575; // @[OneHot.scala 66:30:@37287.4]
  wire [7:0] _T_91640; // @[Mux.scala 19:72:@37311.4]
  wire [15:0] _T_91648; // @[Mux.scala 19:72:@37319.4]
  wire [15:0] _T_91650; // @[Mux.scala 19:72:@37320.4]
  wire [7:0] _T_91657; // @[Mux.scala 19:72:@37327.4]
  wire [15:0] _T_91665; // @[Mux.scala 19:72:@37335.4]
  wire [15:0] _T_91667; // @[Mux.scala 19:72:@37336.4]
  wire [7:0] _T_91674; // @[Mux.scala 19:72:@37343.4]
  wire [15:0] _T_91682; // @[Mux.scala 19:72:@37351.4]
  wire [15:0] _T_91684; // @[Mux.scala 19:72:@37352.4]
  wire [7:0] _T_91691; // @[Mux.scala 19:72:@37359.4]
  wire [15:0] _T_91699; // @[Mux.scala 19:72:@37367.4]
  wire [15:0] _T_91701; // @[Mux.scala 19:72:@37368.4]
  wire [7:0] _T_91708; // @[Mux.scala 19:72:@37375.4]
  wire [15:0] _T_91716; // @[Mux.scala 19:72:@37383.4]
  wire [15:0] _T_91718; // @[Mux.scala 19:72:@37384.4]
  wire [7:0] _T_91725; // @[Mux.scala 19:72:@37391.4]
  wire [15:0] _T_91733; // @[Mux.scala 19:72:@37399.4]
  wire [15:0] _T_91735; // @[Mux.scala 19:72:@37400.4]
  wire [7:0] _T_91742; // @[Mux.scala 19:72:@37407.4]
  wire [15:0] _T_91750; // @[Mux.scala 19:72:@37415.4]
  wire [15:0] _T_91752; // @[Mux.scala 19:72:@37416.4]
  wire [7:0] _T_91759; // @[Mux.scala 19:72:@37423.4]
  wire [15:0] _T_91767; // @[Mux.scala 19:72:@37431.4]
  wire [15:0] _T_91769; // @[Mux.scala 19:72:@37432.4]
  wire [7:0] _T_91776; // @[Mux.scala 19:72:@37439.4]
  wire [15:0] _T_91784; // @[Mux.scala 19:72:@37447.4]
  wire [15:0] _T_91786; // @[Mux.scala 19:72:@37448.4]
  wire [7:0] _T_91793; // @[Mux.scala 19:72:@37455.4]
  wire [15:0] _T_91801; // @[Mux.scala 19:72:@37463.4]
  wire [15:0] _T_91803; // @[Mux.scala 19:72:@37464.4]
  wire [7:0] _T_91810; // @[Mux.scala 19:72:@37471.4]
  wire [15:0] _T_91818; // @[Mux.scala 19:72:@37479.4]
  wire [15:0] _T_91820; // @[Mux.scala 19:72:@37480.4]
  wire [7:0] _T_91827; // @[Mux.scala 19:72:@37487.4]
  wire [15:0] _T_91835; // @[Mux.scala 19:72:@37495.4]
  wire [15:0] _T_91837; // @[Mux.scala 19:72:@37496.4]
  wire [7:0] _T_91844; // @[Mux.scala 19:72:@37503.4]
  wire [15:0] _T_91852; // @[Mux.scala 19:72:@37511.4]
  wire [15:0] _T_91854; // @[Mux.scala 19:72:@37512.4]
  wire [7:0] _T_91861; // @[Mux.scala 19:72:@37519.4]
  wire [15:0] _T_91869; // @[Mux.scala 19:72:@37527.4]
  wire [15:0] _T_91871; // @[Mux.scala 19:72:@37528.4]
  wire [7:0] _T_91878; // @[Mux.scala 19:72:@37535.4]
  wire [15:0] _T_91886; // @[Mux.scala 19:72:@37543.4]
  wire [15:0] _T_91888; // @[Mux.scala 19:72:@37544.4]
  wire [7:0] _T_91895; // @[Mux.scala 19:72:@37551.4]
  wire [15:0] _T_91903; // @[Mux.scala 19:72:@37559.4]
  wire [15:0] _T_91905; // @[Mux.scala 19:72:@37560.4]
  wire [15:0] _T_91906; // @[Mux.scala 19:72:@37561.4]
  wire [15:0] _T_91907; // @[Mux.scala 19:72:@37562.4]
  wire [15:0] _T_91908; // @[Mux.scala 19:72:@37563.4]
  wire [15:0] _T_91909; // @[Mux.scala 19:72:@37564.4]
  wire [15:0] _T_91910; // @[Mux.scala 19:72:@37565.4]
  wire [15:0] _T_91911; // @[Mux.scala 19:72:@37566.4]
  wire [15:0] _T_91912; // @[Mux.scala 19:72:@37567.4]
  wire [15:0] _T_91913; // @[Mux.scala 19:72:@37568.4]
  wire [15:0] _T_91914; // @[Mux.scala 19:72:@37569.4]
  wire [15:0] _T_91915; // @[Mux.scala 19:72:@37570.4]
  wire [15:0] _T_91916; // @[Mux.scala 19:72:@37571.4]
  wire [15:0] _T_91917; // @[Mux.scala 19:72:@37572.4]
  wire [15:0] _T_91918; // @[Mux.scala 19:72:@37573.4]
  wire [15:0] _T_91919; // @[Mux.scala 19:72:@37574.4]
  wire [15:0] _T_91920; // @[Mux.scala 19:72:@37575.4]
  wire  priorityLoadRequest_0; // @[Mux.scala 19:72:@37579.4]
  wire  priorityLoadRequest_1; // @[Mux.scala 19:72:@37581.4]
  wire  priorityLoadRequest_2; // @[Mux.scala 19:72:@37583.4]
  wire  priorityLoadRequest_3; // @[Mux.scala 19:72:@37585.4]
  wire  priorityLoadRequest_4; // @[Mux.scala 19:72:@37587.4]
  wire  priorityLoadRequest_5; // @[Mux.scala 19:72:@37589.4]
  wire  priorityLoadRequest_6; // @[Mux.scala 19:72:@37591.4]
  wire  priorityLoadRequest_7; // @[Mux.scala 19:72:@37593.4]
  wire  priorityLoadRequest_8; // @[Mux.scala 19:72:@37595.4]
  wire  priorityLoadRequest_9; // @[Mux.scala 19:72:@37597.4]
  wire  priorityLoadRequest_10; // @[Mux.scala 19:72:@37599.4]
  wire  priorityLoadRequest_11; // @[Mux.scala 19:72:@37601.4]
  wire  priorityLoadRequest_12; // @[Mux.scala 19:72:@37603.4]
  wire  priorityLoadRequest_13; // @[Mux.scala 19:72:@37605.4]
  wire  priorityLoadRequest_14; // @[Mux.scala 19:72:@37607.4]
  wire  priorityLoadRequest_15; // @[Mux.scala 19:72:@37609.4]
  wire  _GEN_1920; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1921; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1922; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1923; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1924; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1925; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1926; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1927; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1928; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1929; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1930; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1931; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1932; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1933; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1934; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1935; // @[LoadQueue.scala 208:31:@37629.4]
  wire [7:0] _T_92315; // @[LoadQueue.scala 238:58:@37847.8]
  wire [15:0] _T_92323; // @[LoadQueue.scala 238:58:@37855.8]
  wire [7:0] _T_92330; // @[LoadQueue.scala 238:96:@37862.8]
  wire [15:0] _T_92338; // @[LoadQueue.scala 238:96:@37870.8]
  wire  _T_92339; // @[LoadQueue.scala 238:61:@37871.8]
  wire  _T_92340; // @[LoadQueue.scala 237:64:@37872.8]
  wire  _GEN_1969; // @[LoadQueue.scala 230:110:@37804.6]
  wire  bypassRequest_0; // @[LoadQueue.scala 229:71:@37798.4]
  wire  _GEN_1936; // @[LoadQueue.scala 217:34:@37686.6]
  wire  _GEN_1937; // @[LoadQueue.scala 215:23:@37682.4]
  wire [7:0] _T_92399; // @[LoadQueue.scala 238:58:@37929.8]
  wire [15:0] _T_92407; // @[LoadQueue.scala 238:58:@37937.8]
  wire [7:0] _T_92414; // @[LoadQueue.scala 238:96:@37944.8]
  wire [15:0] _T_92422; // @[LoadQueue.scala 238:96:@37952.8]
  wire  _T_92423; // @[LoadQueue.scala 238:61:@37953.8]
  wire  _T_92424; // @[LoadQueue.scala 237:64:@37954.8]
  wire  _GEN_1973; // @[LoadQueue.scala 230:110:@37886.6]
  wire  bypassRequest_1; // @[LoadQueue.scala 229:71:@37880.4]
  wire  _GEN_1938; // @[LoadQueue.scala 217:34:@37693.6]
  wire  _GEN_1939; // @[LoadQueue.scala 215:23:@37689.4]
  wire [7:0] _T_92483; // @[LoadQueue.scala 238:58:@38011.8]
  wire [15:0] _T_92491; // @[LoadQueue.scala 238:58:@38019.8]
  wire [7:0] _T_92498; // @[LoadQueue.scala 238:96:@38026.8]
  wire [15:0] _T_92506; // @[LoadQueue.scala 238:96:@38034.8]
  wire  _T_92507; // @[LoadQueue.scala 238:61:@38035.8]
  wire  _T_92508; // @[LoadQueue.scala 237:64:@38036.8]
  wire  _GEN_1977; // @[LoadQueue.scala 230:110:@37968.6]
  wire  bypassRequest_2; // @[LoadQueue.scala 229:71:@37962.4]
  wire  _GEN_1940; // @[LoadQueue.scala 217:34:@37700.6]
  wire  _GEN_1941; // @[LoadQueue.scala 215:23:@37696.4]
  wire [7:0] _T_92567; // @[LoadQueue.scala 238:58:@38093.8]
  wire [15:0] _T_92575; // @[LoadQueue.scala 238:58:@38101.8]
  wire [7:0] _T_92582; // @[LoadQueue.scala 238:96:@38108.8]
  wire [15:0] _T_92590; // @[LoadQueue.scala 238:96:@38116.8]
  wire  _T_92591; // @[LoadQueue.scala 238:61:@38117.8]
  wire  _T_92592; // @[LoadQueue.scala 237:64:@38118.8]
  wire  _GEN_1981; // @[LoadQueue.scala 230:110:@38050.6]
  wire  bypassRequest_3; // @[LoadQueue.scala 229:71:@38044.4]
  wire  _GEN_1942; // @[LoadQueue.scala 217:34:@37707.6]
  wire  _GEN_1943; // @[LoadQueue.scala 215:23:@37703.4]
  wire [7:0] _T_92651; // @[LoadQueue.scala 238:58:@38175.8]
  wire [15:0] _T_92659; // @[LoadQueue.scala 238:58:@38183.8]
  wire [7:0] _T_92666; // @[LoadQueue.scala 238:96:@38190.8]
  wire [15:0] _T_92674; // @[LoadQueue.scala 238:96:@38198.8]
  wire  _T_92675; // @[LoadQueue.scala 238:61:@38199.8]
  wire  _T_92676; // @[LoadQueue.scala 237:64:@38200.8]
  wire  _GEN_1985; // @[LoadQueue.scala 230:110:@38132.6]
  wire  bypassRequest_4; // @[LoadQueue.scala 229:71:@38126.4]
  wire  _GEN_1944; // @[LoadQueue.scala 217:34:@37714.6]
  wire  _GEN_1945; // @[LoadQueue.scala 215:23:@37710.4]
  wire [7:0] _T_92735; // @[LoadQueue.scala 238:58:@38257.8]
  wire [15:0] _T_92743; // @[LoadQueue.scala 238:58:@38265.8]
  wire [7:0] _T_92750; // @[LoadQueue.scala 238:96:@38272.8]
  wire [15:0] _T_92758; // @[LoadQueue.scala 238:96:@38280.8]
  wire  _T_92759; // @[LoadQueue.scala 238:61:@38281.8]
  wire  _T_92760; // @[LoadQueue.scala 237:64:@38282.8]
  wire  _GEN_1989; // @[LoadQueue.scala 230:110:@38214.6]
  wire  bypassRequest_5; // @[LoadQueue.scala 229:71:@38208.4]
  wire  _GEN_1946; // @[LoadQueue.scala 217:34:@37721.6]
  wire  _GEN_1947; // @[LoadQueue.scala 215:23:@37717.4]
  wire [7:0] _T_92819; // @[LoadQueue.scala 238:58:@38339.8]
  wire [15:0] _T_92827; // @[LoadQueue.scala 238:58:@38347.8]
  wire [7:0] _T_92834; // @[LoadQueue.scala 238:96:@38354.8]
  wire [15:0] _T_92842; // @[LoadQueue.scala 238:96:@38362.8]
  wire  _T_92843; // @[LoadQueue.scala 238:61:@38363.8]
  wire  _T_92844; // @[LoadQueue.scala 237:64:@38364.8]
  wire  _GEN_1993; // @[LoadQueue.scala 230:110:@38296.6]
  wire  bypassRequest_6; // @[LoadQueue.scala 229:71:@38290.4]
  wire  _GEN_1948; // @[LoadQueue.scala 217:34:@37728.6]
  wire  _GEN_1949; // @[LoadQueue.scala 215:23:@37724.4]
  wire [7:0] _T_92903; // @[LoadQueue.scala 238:58:@38421.8]
  wire [15:0] _T_92911; // @[LoadQueue.scala 238:58:@38429.8]
  wire [7:0] _T_92918; // @[LoadQueue.scala 238:96:@38436.8]
  wire [15:0] _T_92926; // @[LoadQueue.scala 238:96:@38444.8]
  wire  _T_92927; // @[LoadQueue.scala 238:61:@38445.8]
  wire  _T_92928; // @[LoadQueue.scala 237:64:@38446.8]
  wire  _GEN_1997; // @[LoadQueue.scala 230:110:@38378.6]
  wire  bypassRequest_7; // @[LoadQueue.scala 229:71:@38372.4]
  wire  _GEN_1950; // @[LoadQueue.scala 217:34:@37735.6]
  wire  _GEN_1951; // @[LoadQueue.scala 215:23:@37731.4]
  wire [7:0] _T_92987; // @[LoadQueue.scala 238:58:@38503.8]
  wire [15:0] _T_92995; // @[LoadQueue.scala 238:58:@38511.8]
  wire [7:0] _T_93002; // @[LoadQueue.scala 238:96:@38518.8]
  wire [15:0] _T_93010; // @[LoadQueue.scala 238:96:@38526.8]
  wire  _T_93011; // @[LoadQueue.scala 238:61:@38527.8]
  wire  _T_93012; // @[LoadQueue.scala 237:64:@38528.8]
  wire  _GEN_2001; // @[LoadQueue.scala 230:110:@38460.6]
  wire  bypassRequest_8; // @[LoadQueue.scala 229:71:@38454.4]
  wire  _GEN_1952; // @[LoadQueue.scala 217:34:@37742.6]
  wire  _GEN_1953; // @[LoadQueue.scala 215:23:@37738.4]
  wire [7:0] _T_93071; // @[LoadQueue.scala 238:58:@38585.8]
  wire [15:0] _T_93079; // @[LoadQueue.scala 238:58:@38593.8]
  wire [7:0] _T_93086; // @[LoadQueue.scala 238:96:@38600.8]
  wire [15:0] _T_93094; // @[LoadQueue.scala 238:96:@38608.8]
  wire  _T_93095; // @[LoadQueue.scala 238:61:@38609.8]
  wire  _T_93096; // @[LoadQueue.scala 237:64:@38610.8]
  wire  _GEN_2005; // @[LoadQueue.scala 230:110:@38542.6]
  wire  bypassRequest_9; // @[LoadQueue.scala 229:71:@38536.4]
  wire  _GEN_1954; // @[LoadQueue.scala 217:34:@37749.6]
  wire  _GEN_1955; // @[LoadQueue.scala 215:23:@37745.4]
  wire [7:0] _T_93155; // @[LoadQueue.scala 238:58:@38667.8]
  wire [15:0] _T_93163; // @[LoadQueue.scala 238:58:@38675.8]
  wire [7:0] _T_93170; // @[LoadQueue.scala 238:96:@38682.8]
  wire [15:0] _T_93178; // @[LoadQueue.scala 238:96:@38690.8]
  wire  _T_93179; // @[LoadQueue.scala 238:61:@38691.8]
  wire  _T_93180; // @[LoadQueue.scala 237:64:@38692.8]
  wire  _GEN_2009; // @[LoadQueue.scala 230:110:@38624.6]
  wire  bypassRequest_10; // @[LoadQueue.scala 229:71:@38618.4]
  wire  _GEN_1956; // @[LoadQueue.scala 217:34:@37756.6]
  wire  _GEN_1957; // @[LoadQueue.scala 215:23:@37752.4]
  wire [7:0] _T_93239; // @[LoadQueue.scala 238:58:@38749.8]
  wire [15:0] _T_93247; // @[LoadQueue.scala 238:58:@38757.8]
  wire [7:0] _T_93254; // @[LoadQueue.scala 238:96:@38764.8]
  wire [15:0] _T_93262; // @[LoadQueue.scala 238:96:@38772.8]
  wire  _T_93263; // @[LoadQueue.scala 238:61:@38773.8]
  wire  _T_93264; // @[LoadQueue.scala 237:64:@38774.8]
  wire  _GEN_2013; // @[LoadQueue.scala 230:110:@38706.6]
  wire  bypassRequest_11; // @[LoadQueue.scala 229:71:@38700.4]
  wire  _GEN_1958; // @[LoadQueue.scala 217:34:@37763.6]
  wire  _GEN_1959; // @[LoadQueue.scala 215:23:@37759.4]
  wire [7:0] _T_93323; // @[LoadQueue.scala 238:58:@38831.8]
  wire [15:0] _T_93331; // @[LoadQueue.scala 238:58:@38839.8]
  wire [7:0] _T_93338; // @[LoadQueue.scala 238:96:@38846.8]
  wire [15:0] _T_93346; // @[LoadQueue.scala 238:96:@38854.8]
  wire  _T_93347; // @[LoadQueue.scala 238:61:@38855.8]
  wire  _T_93348; // @[LoadQueue.scala 237:64:@38856.8]
  wire  _GEN_2017; // @[LoadQueue.scala 230:110:@38788.6]
  wire  bypassRequest_12; // @[LoadQueue.scala 229:71:@38782.4]
  wire  _GEN_1960; // @[LoadQueue.scala 217:34:@37770.6]
  wire  _GEN_1961; // @[LoadQueue.scala 215:23:@37766.4]
  wire [7:0] _T_93407; // @[LoadQueue.scala 238:58:@38913.8]
  wire [15:0] _T_93415; // @[LoadQueue.scala 238:58:@38921.8]
  wire [7:0] _T_93422; // @[LoadQueue.scala 238:96:@38928.8]
  wire [15:0] _T_93430; // @[LoadQueue.scala 238:96:@38936.8]
  wire  _T_93431; // @[LoadQueue.scala 238:61:@38937.8]
  wire  _T_93432; // @[LoadQueue.scala 237:64:@38938.8]
  wire  _GEN_2021; // @[LoadQueue.scala 230:110:@38870.6]
  wire  bypassRequest_13; // @[LoadQueue.scala 229:71:@38864.4]
  wire  _GEN_1962; // @[LoadQueue.scala 217:34:@37777.6]
  wire  _GEN_1963; // @[LoadQueue.scala 215:23:@37773.4]
  wire [7:0] _T_93491; // @[LoadQueue.scala 238:58:@38995.8]
  wire [15:0] _T_93499; // @[LoadQueue.scala 238:58:@39003.8]
  wire [7:0] _T_93506; // @[LoadQueue.scala 238:96:@39010.8]
  wire [15:0] _T_93514; // @[LoadQueue.scala 238:96:@39018.8]
  wire  _T_93515; // @[LoadQueue.scala 238:61:@39019.8]
  wire  _T_93516; // @[LoadQueue.scala 237:64:@39020.8]
  wire  _GEN_2025; // @[LoadQueue.scala 230:110:@38952.6]
  wire  bypassRequest_14; // @[LoadQueue.scala 229:71:@38946.4]
  wire  _GEN_1964; // @[LoadQueue.scala 217:34:@37784.6]
  wire  _GEN_1965; // @[LoadQueue.scala 215:23:@37780.4]
  wire [7:0] _T_93575; // @[LoadQueue.scala 238:58:@39077.8]
  wire [15:0] _T_93583; // @[LoadQueue.scala 238:58:@39085.8]
  wire [7:0] _T_93590; // @[LoadQueue.scala 238:96:@39092.8]
  wire [15:0] _T_93598; // @[LoadQueue.scala 238:96:@39100.8]
  wire  _T_93599; // @[LoadQueue.scala 238:61:@39101.8]
  wire  _T_93600; // @[LoadQueue.scala 237:64:@39102.8]
  wire  _GEN_2029; // @[LoadQueue.scala 230:110:@39034.6]
  wire  bypassRequest_15; // @[LoadQueue.scala 229:71:@39028.4]
  wire  _GEN_1966; // @[LoadQueue.scala 217:34:@37791.6]
  wire  _GEN_1967; // @[LoadQueue.scala 215:23:@37787.4]
  wire  _T_93604; // @[LoadQueue.scala 247:28:@39108.4]
  wire  _T_93605; // @[LoadQueue.scala 247:28:@39109.4]
  wire  _T_93606; // @[LoadQueue.scala 247:28:@39110.4]
  wire  _T_93607; // @[LoadQueue.scala 247:28:@39111.4]
  wire  _T_93608; // @[LoadQueue.scala 247:28:@39112.4]
  wire  _T_93609; // @[LoadQueue.scala 247:28:@39113.4]
  wire  _T_93610; // @[LoadQueue.scala 247:28:@39114.4]
  wire  _T_93611; // @[LoadQueue.scala 247:28:@39115.4]
  wire  _T_93612; // @[LoadQueue.scala 247:28:@39116.4]
  wire  _T_93613; // @[LoadQueue.scala 247:28:@39117.4]
  wire  _T_93614; // @[LoadQueue.scala 247:28:@39118.4]
  wire  _T_93615; // @[LoadQueue.scala 247:28:@39119.4]
  wire  _T_93616; // @[LoadQueue.scala 247:28:@39120.4]
  wire  _T_93617; // @[LoadQueue.scala 247:28:@39121.4]
  wire  _T_93618; // @[LoadQueue.scala 247:28:@39122.4]
  wire [3:0] _T_93635; // @[Mux.scala 31:69:@39124.6]
  wire [3:0] _T_93636; // @[Mux.scala 31:69:@39125.6]
  wire [3:0] _T_93637; // @[Mux.scala 31:69:@39126.6]
  wire [3:0] _T_93638; // @[Mux.scala 31:69:@39127.6]
  wire [3:0] _T_93639; // @[Mux.scala 31:69:@39128.6]
  wire [3:0] _T_93640; // @[Mux.scala 31:69:@39129.6]
  wire [3:0] _T_93641; // @[Mux.scala 31:69:@39130.6]
  wire [3:0] _T_93642; // @[Mux.scala 31:69:@39131.6]
  wire [3:0] _T_93643; // @[Mux.scala 31:69:@39132.6]
  wire [3:0] _T_93644; // @[Mux.scala 31:69:@39133.6]
  wire [3:0] _T_93645; // @[Mux.scala 31:69:@39134.6]
  wire [3:0] _T_93646; // @[Mux.scala 31:69:@39135.6]
  wire [3:0] _T_93647; // @[Mux.scala 31:69:@39136.6]
  wire [3:0] _T_93648; // @[Mux.scala 31:69:@39137.6]
  wire [3:0] _T_93649; // @[Mux.scala 31:69:@39138.6]
  wire [31:0] _GEN_2033; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2034; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2035; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2036; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2037; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2038; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2039; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2040; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2041; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2042; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2043; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2044; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2045; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2046; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2047; // @[LoadQueue.scala 248:24:@39139.6]
  wire  _T_93657; // @[LoadQueue.scala 261:41:@39150.6]
  wire  _GEN_2050; // @[LoadQueue.scala 261:62:@39151.6]
  wire  _GEN_2051; // @[LoadQueue.scala 259:25:@39146.4]
  wire  _T_93660; // @[LoadQueue.scala 261:41:@39158.6]
  wire  _GEN_2052; // @[LoadQueue.scala 261:62:@39159.6]
  wire  _GEN_2053; // @[LoadQueue.scala 259:25:@39154.4]
  wire  _T_93663; // @[LoadQueue.scala 261:41:@39166.6]
  wire  _GEN_2054; // @[LoadQueue.scala 261:62:@39167.6]
  wire  _GEN_2055; // @[LoadQueue.scala 259:25:@39162.4]
  wire  _T_93666; // @[LoadQueue.scala 261:41:@39174.6]
  wire  _GEN_2056; // @[LoadQueue.scala 261:62:@39175.6]
  wire  _GEN_2057; // @[LoadQueue.scala 259:25:@39170.4]
  wire  _T_93669; // @[LoadQueue.scala 261:41:@39182.6]
  wire  _GEN_2058; // @[LoadQueue.scala 261:62:@39183.6]
  wire  _GEN_2059; // @[LoadQueue.scala 259:25:@39178.4]
  wire  _T_93672; // @[LoadQueue.scala 261:41:@39190.6]
  wire  _GEN_2060; // @[LoadQueue.scala 261:62:@39191.6]
  wire  _GEN_2061; // @[LoadQueue.scala 259:25:@39186.4]
  wire  _T_93675; // @[LoadQueue.scala 261:41:@39198.6]
  wire  _GEN_2062; // @[LoadQueue.scala 261:62:@39199.6]
  wire  _GEN_2063; // @[LoadQueue.scala 259:25:@39194.4]
  wire  _T_93678; // @[LoadQueue.scala 261:41:@39206.6]
  wire  _GEN_2064; // @[LoadQueue.scala 261:62:@39207.6]
  wire  _GEN_2065; // @[LoadQueue.scala 259:25:@39202.4]
  wire  _T_93681; // @[LoadQueue.scala 261:41:@39214.6]
  wire  _GEN_2066; // @[LoadQueue.scala 261:62:@39215.6]
  wire  _GEN_2067; // @[LoadQueue.scala 259:25:@39210.4]
  wire  _T_93684; // @[LoadQueue.scala 261:41:@39222.6]
  wire  _GEN_2068; // @[LoadQueue.scala 261:62:@39223.6]
  wire  _GEN_2069; // @[LoadQueue.scala 259:25:@39218.4]
  wire  _T_93687; // @[LoadQueue.scala 261:41:@39230.6]
  wire  _GEN_2070; // @[LoadQueue.scala 261:62:@39231.6]
  wire  _GEN_2071; // @[LoadQueue.scala 259:25:@39226.4]
  wire  _T_93690; // @[LoadQueue.scala 261:41:@39238.6]
  wire  _GEN_2072; // @[LoadQueue.scala 261:62:@39239.6]
  wire  _GEN_2073; // @[LoadQueue.scala 259:25:@39234.4]
  wire  _T_93693; // @[LoadQueue.scala 261:41:@39246.6]
  wire  _GEN_2074; // @[LoadQueue.scala 261:62:@39247.6]
  wire  _GEN_2075; // @[LoadQueue.scala 259:25:@39242.4]
  wire  _T_93696; // @[LoadQueue.scala 261:41:@39254.6]
  wire  _GEN_2076; // @[LoadQueue.scala 261:62:@39255.6]
  wire  _GEN_2077; // @[LoadQueue.scala 259:25:@39250.4]
  wire  _T_93699; // @[LoadQueue.scala 261:41:@39262.6]
  wire  _GEN_2078; // @[LoadQueue.scala 261:62:@39263.6]
  wire  _GEN_2079; // @[LoadQueue.scala 259:25:@39258.4]
  wire  _T_93702; // @[LoadQueue.scala 261:41:@39270.6]
  wire  _GEN_2080; // @[LoadQueue.scala 261:62:@39271.6]
  wire  _GEN_2081; // @[LoadQueue.scala 259:25:@39266.4]
  wire [31:0] _GEN_2082; // @[LoadQueue.scala 269:44:@39278.6]
  wire [31:0] _GEN_2083; // @[LoadQueue.scala 267:32:@39274.4]
  wire [31:0] _GEN_2084; // @[LoadQueue.scala 269:44:@39285.6]
  wire [31:0] _GEN_2085; // @[LoadQueue.scala 267:32:@39281.4]
  wire [31:0] _GEN_2086; // @[LoadQueue.scala 269:44:@39292.6]
  wire [31:0] _GEN_2087; // @[LoadQueue.scala 267:32:@39288.4]
  wire [31:0] _GEN_2088; // @[LoadQueue.scala 269:44:@39299.6]
  wire [31:0] _GEN_2089; // @[LoadQueue.scala 267:32:@39295.4]
  wire [31:0] _GEN_2090; // @[LoadQueue.scala 269:44:@39306.6]
  wire [31:0] _GEN_2091; // @[LoadQueue.scala 267:32:@39302.4]
  wire [31:0] _GEN_2092; // @[LoadQueue.scala 269:44:@39313.6]
  wire [31:0] _GEN_2093; // @[LoadQueue.scala 267:32:@39309.4]
  wire [31:0] _GEN_2094; // @[LoadQueue.scala 269:44:@39320.6]
  wire [31:0] _GEN_2095; // @[LoadQueue.scala 267:32:@39316.4]
  wire [31:0] _GEN_2096; // @[LoadQueue.scala 269:44:@39327.6]
  wire [31:0] _GEN_2097; // @[LoadQueue.scala 267:32:@39323.4]
  wire [31:0] _GEN_2098; // @[LoadQueue.scala 269:44:@39334.6]
  wire [31:0] _GEN_2099; // @[LoadQueue.scala 267:32:@39330.4]
  wire [31:0] _GEN_2100; // @[LoadQueue.scala 269:44:@39341.6]
  wire [31:0] _GEN_2101; // @[LoadQueue.scala 267:32:@39337.4]
  wire [31:0] _GEN_2102; // @[LoadQueue.scala 269:44:@39348.6]
  wire [31:0] _GEN_2103; // @[LoadQueue.scala 267:32:@39344.4]
  wire [31:0] _GEN_2104; // @[LoadQueue.scala 269:44:@39355.6]
  wire [31:0] _GEN_2105; // @[LoadQueue.scala 267:32:@39351.4]
  wire [31:0] _GEN_2106; // @[LoadQueue.scala 269:44:@39362.6]
  wire [31:0] _GEN_2107; // @[LoadQueue.scala 267:32:@39358.4]
  wire [31:0] _GEN_2108; // @[LoadQueue.scala 269:44:@39369.6]
  wire [31:0] _GEN_2109; // @[LoadQueue.scala 267:32:@39365.4]
  wire [31:0] _GEN_2110; // @[LoadQueue.scala 269:44:@39376.6]
  wire [31:0] _GEN_2111; // @[LoadQueue.scala 267:32:@39372.4]
  wire [31:0] _GEN_2112; // @[LoadQueue.scala 269:44:@39383.6]
  wire [31:0] _GEN_2113; // @[LoadQueue.scala 267:32:@39379.4]
  wire  entriesPorts_0_0; // @[LoadQueue.scala 286:69:@39387.4]
  wire  entriesPorts_0_1; // @[LoadQueue.scala 286:69:@39389.4]
  wire  entriesPorts_0_2; // @[LoadQueue.scala 286:69:@39391.4]
  wire  entriesPorts_0_3; // @[LoadQueue.scala 286:69:@39393.4]
  wire  entriesPorts_0_4; // @[LoadQueue.scala 286:69:@39395.4]
  wire  entriesPorts_0_5; // @[LoadQueue.scala 286:69:@39397.4]
  wire  entriesPorts_0_6; // @[LoadQueue.scala 286:69:@39399.4]
  wire  entriesPorts_0_7; // @[LoadQueue.scala 286:69:@39401.4]
  wire  entriesPorts_0_8; // @[LoadQueue.scala 286:69:@39403.4]
  wire  entriesPorts_0_9; // @[LoadQueue.scala 286:69:@39405.4]
  wire  entriesPorts_0_10; // @[LoadQueue.scala 286:69:@39407.4]
  wire  entriesPorts_0_11; // @[LoadQueue.scala 286:69:@39409.4]
  wire  entriesPorts_0_12; // @[LoadQueue.scala 286:69:@39411.4]
  wire  entriesPorts_0_13; // @[LoadQueue.scala 286:69:@39413.4]
  wire  entriesPorts_0_14; // @[LoadQueue.scala 286:69:@39415.4]
  wire  entriesPorts_0_15; // @[LoadQueue.scala 286:69:@39417.4]
  wire  _T_94435; // @[LoadQueue.scala 298:86:@39453.4]
  wire  _T_94436; // @[LoadQueue.scala 298:83:@39454.4]
  wire  _T_94438; // @[LoadQueue.scala 298:86:@39455.4]
  wire  _T_94439; // @[LoadQueue.scala 298:83:@39456.4]
  wire  _T_94441; // @[LoadQueue.scala 298:86:@39457.4]
  wire  _T_94442; // @[LoadQueue.scala 298:83:@39458.4]
  wire  _T_94444; // @[LoadQueue.scala 298:86:@39459.4]
  wire  _T_94445; // @[LoadQueue.scala 298:83:@39460.4]
  wire  _T_94447; // @[LoadQueue.scala 298:86:@39461.4]
  wire  _T_94448; // @[LoadQueue.scala 298:83:@39462.4]
  wire  _T_94450; // @[LoadQueue.scala 298:86:@39463.4]
  wire  _T_94451; // @[LoadQueue.scala 298:83:@39464.4]
  wire  _T_94453; // @[LoadQueue.scala 298:86:@39465.4]
  wire  _T_94454; // @[LoadQueue.scala 298:83:@39466.4]
  wire  _T_94456; // @[LoadQueue.scala 298:86:@39467.4]
  wire  _T_94457; // @[LoadQueue.scala 298:83:@39468.4]
  wire  _T_94459; // @[LoadQueue.scala 298:86:@39469.4]
  wire  _T_94460; // @[LoadQueue.scala 298:83:@39470.4]
  wire  _T_94462; // @[LoadQueue.scala 298:86:@39471.4]
  wire  _T_94463; // @[LoadQueue.scala 298:83:@39472.4]
  wire  _T_94465; // @[LoadQueue.scala 298:86:@39473.4]
  wire  _T_94466; // @[LoadQueue.scala 298:83:@39474.4]
  wire  _T_94468; // @[LoadQueue.scala 298:86:@39475.4]
  wire  _T_94469; // @[LoadQueue.scala 298:83:@39476.4]
  wire  _T_94471; // @[LoadQueue.scala 298:86:@39477.4]
  wire  _T_94472; // @[LoadQueue.scala 298:83:@39478.4]
  wire  _T_94474; // @[LoadQueue.scala 298:86:@39479.4]
  wire  _T_94475; // @[LoadQueue.scala 298:83:@39480.4]
  wire  _T_94477; // @[LoadQueue.scala 298:86:@39481.4]
  wire  _T_94478; // @[LoadQueue.scala 298:83:@39482.4]
  wire  _T_94480; // @[LoadQueue.scala 298:86:@39483.4]
  wire  _T_94481; // @[LoadQueue.scala 298:83:@39484.4]
  wire [15:0] _T_94564; // @[Mux.scala 31:69:@39538.4]
  wire [15:0] _T_94565; // @[Mux.scala 31:69:@39539.4]
  wire [15:0] _T_94566; // @[Mux.scala 31:69:@39540.4]
  wire [15:0] _T_94567; // @[Mux.scala 31:69:@39541.4]
  wire [15:0] _T_94568; // @[Mux.scala 31:69:@39542.4]
  wire [15:0] _T_94569; // @[Mux.scala 31:69:@39543.4]
  wire [15:0] _T_94570; // @[Mux.scala 31:69:@39544.4]
  wire [15:0] _T_94571; // @[Mux.scala 31:69:@39545.4]
  wire [15:0] _T_94572; // @[Mux.scala 31:69:@39546.4]
  wire [15:0] _T_94573; // @[Mux.scala 31:69:@39547.4]
  wire [15:0] _T_94574; // @[Mux.scala 31:69:@39548.4]
  wire [15:0] _T_94575; // @[Mux.scala 31:69:@39549.4]
  wire [15:0] _T_94576; // @[Mux.scala 31:69:@39550.4]
  wire [15:0] _T_94577; // @[Mux.scala 31:69:@39551.4]
  wire [15:0] _T_94578; // @[Mux.scala 31:69:@39552.4]
  wire [15:0] _T_94579; // @[Mux.scala 31:69:@39553.4]
  wire  _T_94580; // @[OneHot.scala 66:30:@39554.4]
  wire  _T_94581; // @[OneHot.scala 66:30:@39555.4]
  wire  _T_94582; // @[OneHot.scala 66:30:@39556.4]
  wire  _T_94583; // @[OneHot.scala 66:30:@39557.4]
  wire  _T_94584; // @[OneHot.scala 66:30:@39558.4]
  wire  _T_94585; // @[OneHot.scala 66:30:@39559.4]
  wire  _T_94586; // @[OneHot.scala 66:30:@39560.4]
  wire  _T_94587; // @[OneHot.scala 66:30:@39561.4]
  wire  _T_94588; // @[OneHot.scala 66:30:@39562.4]
  wire  _T_94589; // @[OneHot.scala 66:30:@39563.4]
  wire  _T_94590; // @[OneHot.scala 66:30:@39564.4]
  wire  _T_94591; // @[OneHot.scala 66:30:@39565.4]
  wire  _T_94592; // @[OneHot.scala 66:30:@39566.4]
  wire  _T_94593; // @[OneHot.scala 66:30:@39567.4]
  wire  _T_94594; // @[OneHot.scala 66:30:@39568.4]
  wire  _T_94595; // @[OneHot.scala 66:30:@39569.4]
  wire [15:0] _T_94636; // @[Mux.scala 31:69:@39587.4]
  wire [15:0] _T_94637; // @[Mux.scala 31:69:@39588.4]
  wire [15:0] _T_94638; // @[Mux.scala 31:69:@39589.4]
  wire [15:0] _T_94639; // @[Mux.scala 31:69:@39590.4]
  wire [15:0] _T_94640; // @[Mux.scala 31:69:@39591.4]
  wire [15:0] _T_94641; // @[Mux.scala 31:69:@39592.4]
  wire [15:0] _T_94642; // @[Mux.scala 31:69:@39593.4]
  wire [15:0] _T_94643; // @[Mux.scala 31:69:@39594.4]
  wire [15:0] _T_94644; // @[Mux.scala 31:69:@39595.4]
  wire [15:0] _T_94645; // @[Mux.scala 31:69:@39596.4]
  wire [15:0] _T_94646; // @[Mux.scala 31:69:@39597.4]
  wire [15:0] _T_94647; // @[Mux.scala 31:69:@39598.4]
  wire [15:0] _T_94648; // @[Mux.scala 31:69:@39599.4]
  wire [15:0] _T_94649; // @[Mux.scala 31:69:@39600.4]
  wire [15:0] _T_94650; // @[Mux.scala 31:69:@39601.4]
  wire [15:0] _T_94651; // @[Mux.scala 31:69:@39602.4]
  wire  _T_94652; // @[OneHot.scala 66:30:@39603.4]
  wire  _T_94653; // @[OneHot.scala 66:30:@39604.4]
  wire  _T_94654; // @[OneHot.scala 66:30:@39605.4]
  wire  _T_94655; // @[OneHot.scala 66:30:@39606.4]
  wire  _T_94656; // @[OneHot.scala 66:30:@39607.4]
  wire  _T_94657; // @[OneHot.scala 66:30:@39608.4]
  wire  _T_94658; // @[OneHot.scala 66:30:@39609.4]
  wire  _T_94659; // @[OneHot.scala 66:30:@39610.4]
  wire  _T_94660; // @[OneHot.scala 66:30:@39611.4]
  wire  _T_94661; // @[OneHot.scala 66:30:@39612.4]
  wire  _T_94662; // @[OneHot.scala 66:30:@39613.4]
  wire  _T_94663; // @[OneHot.scala 66:30:@39614.4]
  wire  _T_94664; // @[OneHot.scala 66:30:@39615.4]
  wire  _T_94665; // @[OneHot.scala 66:30:@39616.4]
  wire  _T_94666; // @[OneHot.scala 66:30:@39617.4]
  wire  _T_94667; // @[OneHot.scala 66:30:@39618.4]
  wire [15:0] _T_94708; // @[Mux.scala 31:69:@39636.4]
  wire [15:0] _T_94709; // @[Mux.scala 31:69:@39637.4]
  wire [15:0] _T_94710; // @[Mux.scala 31:69:@39638.4]
  wire [15:0] _T_94711; // @[Mux.scala 31:69:@39639.4]
  wire [15:0] _T_94712; // @[Mux.scala 31:69:@39640.4]
  wire [15:0] _T_94713; // @[Mux.scala 31:69:@39641.4]
  wire [15:0] _T_94714; // @[Mux.scala 31:69:@39642.4]
  wire [15:0] _T_94715; // @[Mux.scala 31:69:@39643.4]
  wire [15:0] _T_94716; // @[Mux.scala 31:69:@39644.4]
  wire [15:0] _T_94717; // @[Mux.scala 31:69:@39645.4]
  wire [15:0] _T_94718; // @[Mux.scala 31:69:@39646.4]
  wire [15:0] _T_94719; // @[Mux.scala 31:69:@39647.4]
  wire [15:0] _T_94720; // @[Mux.scala 31:69:@39648.4]
  wire [15:0] _T_94721; // @[Mux.scala 31:69:@39649.4]
  wire [15:0] _T_94722; // @[Mux.scala 31:69:@39650.4]
  wire [15:0] _T_94723; // @[Mux.scala 31:69:@39651.4]
  wire  _T_94724; // @[OneHot.scala 66:30:@39652.4]
  wire  _T_94725; // @[OneHot.scala 66:30:@39653.4]
  wire  _T_94726; // @[OneHot.scala 66:30:@39654.4]
  wire  _T_94727; // @[OneHot.scala 66:30:@39655.4]
  wire  _T_94728; // @[OneHot.scala 66:30:@39656.4]
  wire  _T_94729; // @[OneHot.scala 66:30:@39657.4]
  wire  _T_94730; // @[OneHot.scala 66:30:@39658.4]
  wire  _T_94731; // @[OneHot.scala 66:30:@39659.4]
  wire  _T_94732; // @[OneHot.scala 66:30:@39660.4]
  wire  _T_94733; // @[OneHot.scala 66:30:@39661.4]
  wire  _T_94734; // @[OneHot.scala 66:30:@39662.4]
  wire  _T_94735; // @[OneHot.scala 66:30:@39663.4]
  wire  _T_94736; // @[OneHot.scala 66:30:@39664.4]
  wire  _T_94737; // @[OneHot.scala 66:30:@39665.4]
  wire  _T_94738; // @[OneHot.scala 66:30:@39666.4]
  wire  _T_94739; // @[OneHot.scala 66:30:@39667.4]
  wire [15:0] _T_94780; // @[Mux.scala 31:69:@39685.4]
  wire [15:0] _T_94781; // @[Mux.scala 31:69:@39686.4]
  wire [15:0] _T_94782; // @[Mux.scala 31:69:@39687.4]
  wire [15:0] _T_94783; // @[Mux.scala 31:69:@39688.4]
  wire [15:0] _T_94784; // @[Mux.scala 31:69:@39689.4]
  wire [15:0] _T_94785; // @[Mux.scala 31:69:@39690.4]
  wire [15:0] _T_94786; // @[Mux.scala 31:69:@39691.4]
  wire [15:0] _T_94787; // @[Mux.scala 31:69:@39692.4]
  wire [15:0] _T_94788; // @[Mux.scala 31:69:@39693.4]
  wire [15:0] _T_94789; // @[Mux.scala 31:69:@39694.4]
  wire [15:0] _T_94790; // @[Mux.scala 31:69:@39695.4]
  wire [15:0] _T_94791; // @[Mux.scala 31:69:@39696.4]
  wire [15:0] _T_94792; // @[Mux.scala 31:69:@39697.4]
  wire [15:0] _T_94793; // @[Mux.scala 31:69:@39698.4]
  wire [15:0] _T_94794; // @[Mux.scala 31:69:@39699.4]
  wire [15:0] _T_94795; // @[Mux.scala 31:69:@39700.4]
  wire  _T_94796; // @[OneHot.scala 66:30:@39701.4]
  wire  _T_94797; // @[OneHot.scala 66:30:@39702.4]
  wire  _T_94798; // @[OneHot.scala 66:30:@39703.4]
  wire  _T_94799; // @[OneHot.scala 66:30:@39704.4]
  wire  _T_94800; // @[OneHot.scala 66:30:@39705.4]
  wire  _T_94801; // @[OneHot.scala 66:30:@39706.4]
  wire  _T_94802; // @[OneHot.scala 66:30:@39707.4]
  wire  _T_94803; // @[OneHot.scala 66:30:@39708.4]
  wire  _T_94804; // @[OneHot.scala 66:30:@39709.4]
  wire  _T_94805; // @[OneHot.scala 66:30:@39710.4]
  wire  _T_94806; // @[OneHot.scala 66:30:@39711.4]
  wire  _T_94807; // @[OneHot.scala 66:30:@39712.4]
  wire  _T_94808; // @[OneHot.scala 66:30:@39713.4]
  wire  _T_94809; // @[OneHot.scala 66:30:@39714.4]
  wire  _T_94810; // @[OneHot.scala 66:30:@39715.4]
  wire  _T_94811; // @[OneHot.scala 66:30:@39716.4]
  wire [15:0] _T_94852; // @[Mux.scala 31:69:@39734.4]
  wire [15:0] _T_94853; // @[Mux.scala 31:69:@39735.4]
  wire [15:0] _T_94854; // @[Mux.scala 31:69:@39736.4]
  wire [15:0] _T_94855; // @[Mux.scala 31:69:@39737.4]
  wire [15:0] _T_94856; // @[Mux.scala 31:69:@39738.4]
  wire [15:0] _T_94857; // @[Mux.scala 31:69:@39739.4]
  wire [15:0] _T_94858; // @[Mux.scala 31:69:@39740.4]
  wire [15:0] _T_94859; // @[Mux.scala 31:69:@39741.4]
  wire [15:0] _T_94860; // @[Mux.scala 31:69:@39742.4]
  wire [15:0] _T_94861; // @[Mux.scala 31:69:@39743.4]
  wire [15:0] _T_94862; // @[Mux.scala 31:69:@39744.4]
  wire [15:0] _T_94863; // @[Mux.scala 31:69:@39745.4]
  wire [15:0] _T_94864; // @[Mux.scala 31:69:@39746.4]
  wire [15:0] _T_94865; // @[Mux.scala 31:69:@39747.4]
  wire [15:0] _T_94866; // @[Mux.scala 31:69:@39748.4]
  wire [15:0] _T_94867; // @[Mux.scala 31:69:@39749.4]
  wire  _T_94868; // @[OneHot.scala 66:30:@39750.4]
  wire  _T_94869; // @[OneHot.scala 66:30:@39751.4]
  wire  _T_94870; // @[OneHot.scala 66:30:@39752.4]
  wire  _T_94871; // @[OneHot.scala 66:30:@39753.4]
  wire  _T_94872; // @[OneHot.scala 66:30:@39754.4]
  wire  _T_94873; // @[OneHot.scala 66:30:@39755.4]
  wire  _T_94874; // @[OneHot.scala 66:30:@39756.4]
  wire  _T_94875; // @[OneHot.scala 66:30:@39757.4]
  wire  _T_94876; // @[OneHot.scala 66:30:@39758.4]
  wire  _T_94877; // @[OneHot.scala 66:30:@39759.4]
  wire  _T_94878; // @[OneHot.scala 66:30:@39760.4]
  wire  _T_94879; // @[OneHot.scala 66:30:@39761.4]
  wire  _T_94880; // @[OneHot.scala 66:30:@39762.4]
  wire  _T_94881; // @[OneHot.scala 66:30:@39763.4]
  wire  _T_94882; // @[OneHot.scala 66:30:@39764.4]
  wire  _T_94883; // @[OneHot.scala 66:30:@39765.4]
  wire [15:0] _T_94924; // @[Mux.scala 31:69:@39783.4]
  wire [15:0] _T_94925; // @[Mux.scala 31:69:@39784.4]
  wire [15:0] _T_94926; // @[Mux.scala 31:69:@39785.4]
  wire [15:0] _T_94927; // @[Mux.scala 31:69:@39786.4]
  wire [15:0] _T_94928; // @[Mux.scala 31:69:@39787.4]
  wire [15:0] _T_94929; // @[Mux.scala 31:69:@39788.4]
  wire [15:0] _T_94930; // @[Mux.scala 31:69:@39789.4]
  wire [15:0] _T_94931; // @[Mux.scala 31:69:@39790.4]
  wire [15:0] _T_94932; // @[Mux.scala 31:69:@39791.4]
  wire [15:0] _T_94933; // @[Mux.scala 31:69:@39792.4]
  wire [15:0] _T_94934; // @[Mux.scala 31:69:@39793.4]
  wire [15:0] _T_94935; // @[Mux.scala 31:69:@39794.4]
  wire [15:0] _T_94936; // @[Mux.scala 31:69:@39795.4]
  wire [15:0] _T_94937; // @[Mux.scala 31:69:@39796.4]
  wire [15:0] _T_94938; // @[Mux.scala 31:69:@39797.4]
  wire [15:0] _T_94939; // @[Mux.scala 31:69:@39798.4]
  wire  _T_94940; // @[OneHot.scala 66:30:@39799.4]
  wire  _T_94941; // @[OneHot.scala 66:30:@39800.4]
  wire  _T_94942; // @[OneHot.scala 66:30:@39801.4]
  wire  _T_94943; // @[OneHot.scala 66:30:@39802.4]
  wire  _T_94944; // @[OneHot.scala 66:30:@39803.4]
  wire  _T_94945; // @[OneHot.scala 66:30:@39804.4]
  wire  _T_94946; // @[OneHot.scala 66:30:@39805.4]
  wire  _T_94947; // @[OneHot.scala 66:30:@39806.4]
  wire  _T_94948; // @[OneHot.scala 66:30:@39807.4]
  wire  _T_94949; // @[OneHot.scala 66:30:@39808.4]
  wire  _T_94950; // @[OneHot.scala 66:30:@39809.4]
  wire  _T_94951; // @[OneHot.scala 66:30:@39810.4]
  wire  _T_94952; // @[OneHot.scala 66:30:@39811.4]
  wire  _T_94953; // @[OneHot.scala 66:30:@39812.4]
  wire  _T_94954; // @[OneHot.scala 66:30:@39813.4]
  wire  _T_94955; // @[OneHot.scala 66:30:@39814.4]
  wire [15:0] _T_94996; // @[Mux.scala 31:69:@39832.4]
  wire [15:0] _T_94997; // @[Mux.scala 31:69:@39833.4]
  wire [15:0] _T_94998; // @[Mux.scala 31:69:@39834.4]
  wire [15:0] _T_94999; // @[Mux.scala 31:69:@39835.4]
  wire [15:0] _T_95000; // @[Mux.scala 31:69:@39836.4]
  wire [15:0] _T_95001; // @[Mux.scala 31:69:@39837.4]
  wire [15:0] _T_95002; // @[Mux.scala 31:69:@39838.4]
  wire [15:0] _T_95003; // @[Mux.scala 31:69:@39839.4]
  wire [15:0] _T_95004; // @[Mux.scala 31:69:@39840.4]
  wire [15:0] _T_95005; // @[Mux.scala 31:69:@39841.4]
  wire [15:0] _T_95006; // @[Mux.scala 31:69:@39842.4]
  wire [15:0] _T_95007; // @[Mux.scala 31:69:@39843.4]
  wire [15:0] _T_95008; // @[Mux.scala 31:69:@39844.4]
  wire [15:0] _T_95009; // @[Mux.scala 31:69:@39845.4]
  wire [15:0] _T_95010; // @[Mux.scala 31:69:@39846.4]
  wire [15:0] _T_95011; // @[Mux.scala 31:69:@39847.4]
  wire  _T_95012; // @[OneHot.scala 66:30:@39848.4]
  wire  _T_95013; // @[OneHot.scala 66:30:@39849.4]
  wire  _T_95014; // @[OneHot.scala 66:30:@39850.4]
  wire  _T_95015; // @[OneHot.scala 66:30:@39851.4]
  wire  _T_95016; // @[OneHot.scala 66:30:@39852.4]
  wire  _T_95017; // @[OneHot.scala 66:30:@39853.4]
  wire  _T_95018; // @[OneHot.scala 66:30:@39854.4]
  wire  _T_95019; // @[OneHot.scala 66:30:@39855.4]
  wire  _T_95020; // @[OneHot.scala 66:30:@39856.4]
  wire  _T_95021; // @[OneHot.scala 66:30:@39857.4]
  wire  _T_95022; // @[OneHot.scala 66:30:@39858.4]
  wire  _T_95023; // @[OneHot.scala 66:30:@39859.4]
  wire  _T_95024; // @[OneHot.scala 66:30:@39860.4]
  wire  _T_95025; // @[OneHot.scala 66:30:@39861.4]
  wire  _T_95026; // @[OneHot.scala 66:30:@39862.4]
  wire  _T_95027; // @[OneHot.scala 66:30:@39863.4]
  wire [15:0] _T_95068; // @[Mux.scala 31:69:@39881.4]
  wire [15:0] _T_95069; // @[Mux.scala 31:69:@39882.4]
  wire [15:0] _T_95070; // @[Mux.scala 31:69:@39883.4]
  wire [15:0] _T_95071; // @[Mux.scala 31:69:@39884.4]
  wire [15:0] _T_95072; // @[Mux.scala 31:69:@39885.4]
  wire [15:0] _T_95073; // @[Mux.scala 31:69:@39886.4]
  wire [15:0] _T_95074; // @[Mux.scala 31:69:@39887.4]
  wire [15:0] _T_95075; // @[Mux.scala 31:69:@39888.4]
  wire [15:0] _T_95076; // @[Mux.scala 31:69:@39889.4]
  wire [15:0] _T_95077; // @[Mux.scala 31:69:@39890.4]
  wire [15:0] _T_95078; // @[Mux.scala 31:69:@39891.4]
  wire [15:0] _T_95079; // @[Mux.scala 31:69:@39892.4]
  wire [15:0] _T_95080; // @[Mux.scala 31:69:@39893.4]
  wire [15:0] _T_95081; // @[Mux.scala 31:69:@39894.4]
  wire [15:0] _T_95082; // @[Mux.scala 31:69:@39895.4]
  wire [15:0] _T_95083; // @[Mux.scala 31:69:@39896.4]
  wire  _T_95084; // @[OneHot.scala 66:30:@39897.4]
  wire  _T_95085; // @[OneHot.scala 66:30:@39898.4]
  wire  _T_95086; // @[OneHot.scala 66:30:@39899.4]
  wire  _T_95087; // @[OneHot.scala 66:30:@39900.4]
  wire  _T_95088; // @[OneHot.scala 66:30:@39901.4]
  wire  _T_95089; // @[OneHot.scala 66:30:@39902.4]
  wire  _T_95090; // @[OneHot.scala 66:30:@39903.4]
  wire  _T_95091; // @[OneHot.scala 66:30:@39904.4]
  wire  _T_95092; // @[OneHot.scala 66:30:@39905.4]
  wire  _T_95093; // @[OneHot.scala 66:30:@39906.4]
  wire  _T_95094; // @[OneHot.scala 66:30:@39907.4]
  wire  _T_95095; // @[OneHot.scala 66:30:@39908.4]
  wire  _T_95096; // @[OneHot.scala 66:30:@39909.4]
  wire  _T_95097; // @[OneHot.scala 66:30:@39910.4]
  wire  _T_95098; // @[OneHot.scala 66:30:@39911.4]
  wire  _T_95099; // @[OneHot.scala 66:30:@39912.4]
  wire [15:0] _T_95140; // @[Mux.scala 31:69:@39930.4]
  wire [15:0] _T_95141; // @[Mux.scala 31:69:@39931.4]
  wire [15:0] _T_95142; // @[Mux.scala 31:69:@39932.4]
  wire [15:0] _T_95143; // @[Mux.scala 31:69:@39933.4]
  wire [15:0] _T_95144; // @[Mux.scala 31:69:@39934.4]
  wire [15:0] _T_95145; // @[Mux.scala 31:69:@39935.4]
  wire [15:0] _T_95146; // @[Mux.scala 31:69:@39936.4]
  wire [15:0] _T_95147; // @[Mux.scala 31:69:@39937.4]
  wire [15:0] _T_95148; // @[Mux.scala 31:69:@39938.4]
  wire [15:0] _T_95149; // @[Mux.scala 31:69:@39939.4]
  wire [15:0] _T_95150; // @[Mux.scala 31:69:@39940.4]
  wire [15:0] _T_95151; // @[Mux.scala 31:69:@39941.4]
  wire [15:0] _T_95152; // @[Mux.scala 31:69:@39942.4]
  wire [15:0] _T_95153; // @[Mux.scala 31:69:@39943.4]
  wire [15:0] _T_95154; // @[Mux.scala 31:69:@39944.4]
  wire [15:0] _T_95155; // @[Mux.scala 31:69:@39945.4]
  wire  _T_95156; // @[OneHot.scala 66:30:@39946.4]
  wire  _T_95157; // @[OneHot.scala 66:30:@39947.4]
  wire  _T_95158; // @[OneHot.scala 66:30:@39948.4]
  wire  _T_95159; // @[OneHot.scala 66:30:@39949.4]
  wire  _T_95160; // @[OneHot.scala 66:30:@39950.4]
  wire  _T_95161; // @[OneHot.scala 66:30:@39951.4]
  wire  _T_95162; // @[OneHot.scala 66:30:@39952.4]
  wire  _T_95163; // @[OneHot.scala 66:30:@39953.4]
  wire  _T_95164; // @[OneHot.scala 66:30:@39954.4]
  wire  _T_95165; // @[OneHot.scala 66:30:@39955.4]
  wire  _T_95166; // @[OneHot.scala 66:30:@39956.4]
  wire  _T_95167; // @[OneHot.scala 66:30:@39957.4]
  wire  _T_95168; // @[OneHot.scala 66:30:@39958.4]
  wire  _T_95169; // @[OneHot.scala 66:30:@39959.4]
  wire  _T_95170; // @[OneHot.scala 66:30:@39960.4]
  wire  _T_95171; // @[OneHot.scala 66:30:@39961.4]
  wire [15:0] _T_95212; // @[Mux.scala 31:69:@39979.4]
  wire [15:0] _T_95213; // @[Mux.scala 31:69:@39980.4]
  wire [15:0] _T_95214; // @[Mux.scala 31:69:@39981.4]
  wire [15:0] _T_95215; // @[Mux.scala 31:69:@39982.4]
  wire [15:0] _T_95216; // @[Mux.scala 31:69:@39983.4]
  wire [15:0] _T_95217; // @[Mux.scala 31:69:@39984.4]
  wire [15:0] _T_95218; // @[Mux.scala 31:69:@39985.4]
  wire [15:0] _T_95219; // @[Mux.scala 31:69:@39986.4]
  wire [15:0] _T_95220; // @[Mux.scala 31:69:@39987.4]
  wire [15:0] _T_95221; // @[Mux.scala 31:69:@39988.4]
  wire [15:0] _T_95222; // @[Mux.scala 31:69:@39989.4]
  wire [15:0] _T_95223; // @[Mux.scala 31:69:@39990.4]
  wire [15:0] _T_95224; // @[Mux.scala 31:69:@39991.4]
  wire [15:0] _T_95225; // @[Mux.scala 31:69:@39992.4]
  wire [15:0] _T_95226; // @[Mux.scala 31:69:@39993.4]
  wire [15:0] _T_95227; // @[Mux.scala 31:69:@39994.4]
  wire  _T_95228; // @[OneHot.scala 66:30:@39995.4]
  wire  _T_95229; // @[OneHot.scala 66:30:@39996.4]
  wire  _T_95230; // @[OneHot.scala 66:30:@39997.4]
  wire  _T_95231; // @[OneHot.scala 66:30:@39998.4]
  wire  _T_95232; // @[OneHot.scala 66:30:@39999.4]
  wire  _T_95233; // @[OneHot.scala 66:30:@40000.4]
  wire  _T_95234; // @[OneHot.scala 66:30:@40001.4]
  wire  _T_95235; // @[OneHot.scala 66:30:@40002.4]
  wire  _T_95236; // @[OneHot.scala 66:30:@40003.4]
  wire  _T_95237; // @[OneHot.scala 66:30:@40004.4]
  wire  _T_95238; // @[OneHot.scala 66:30:@40005.4]
  wire  _T_95239; // @[OneHot.scala 66:30:@40006.4]
  wire  _T_95240; // @[OneHot.scala 66:30:@40007.4]
  wire  _T_95241; // @[OneHot.scala 66:30:@40008.4]
  wire  _T_95242; // @[OneHot.scala 66:30:@40009.4]
  wire  _T_95243; // @[OneHot.scala 66:30:@40010.4]
  wire [15:0] _T_95284; // @[Mux.scala 31:69:@40028.4]
  wire [15:0] _T_95285; // @[Mux.scala 31:69:@40029.4]
  wire [15:0] _T_95286; // @[Mux.scala 31:69:@40030.4]
  wire [15:0] _T_95287; // @[Mux.scala 31:69:@40031.4]
  wire [15:0] _T_95288; // @[Mux.scala 31:69:@40032.4]
  wire [15:0] _T_95289; // @[Mux.scala 31:69:@40033.4]
  wire [15:0] _T_95290; // @[Mux.scala 31:69:@40034.4]
  wire [15:0] _T_95291; // @[Mux.scala 31:69:@40035.4]
  wire [15:0] _T_95292; // @[Mux.scala 31:69:@40036.4]
  wire [15:0] _T_95293; // @[Mux.scala 31:69:@40037.4]
  wire [15:0] _T_95294; // @[Mux.scala 31:69:@40038.4]
  wire [15:0] _T_95295; // @[Mux.scala 31:69:@40039.4]
  wire [15:0] _T_95296; // @[Mux.scala 31:69:@40040.4]
  wire [15:0] _T_95297; // @[Mux.scala 31:69:@40041.4]
  wire [15:0] _T_95298; // @[Mux.scala 31:69:@40042.4]
  wire [15:0] _T_95299; // @[Mux.scala 31:69:@40043.4]
  wire  _T_95300; // @[OneHot.scala 66:30:@40044.4]
  wire  _T_95301; // @[OneHot.scala 66:30:@40045.4]
  wire  _T_95302; // @[OneHot.scala 66:30:@40046.4]
  wire  _T_95303; // @[OneHot.scala 66:30:@40047.4]
  wire  _T_95304; // @[OneHot.scala 66:30:@40048.4]
  wire  _T_95305; // @[OneHot.scala 66:30:@40049.4]
  wire  _T_95306; // @[OneHot.scala 66:30:@40050.4]
  wire  _T_95307; // @[OneHot.scala 66:30:@40051.4]
  wire  _T_95308; // @[OneHot.scala 66:30:@40052.4]
  wire  _T_95309; // @[OneHot.scala 66:30:@40053.4]
  wire  _T_95310; // @[OneHot.scala 66:30:@40054.4]
  wire  _T_95311; // @[OneHot.scala 66:30:@40055.4]
  wire  _T_95312; // @[OneHot.scala 66:30:@40056.4]
  wire  _T_95313; // @[OneHot.scala 66:30:@40057.4]
  wire  _T_95314; // @[OneHot.scala 66:30:@40058.4]
  wire  _T_95315; // @[OneHot.scala 66:30:@40059.4]
  wire [15:0] _T_95356; // @[Mux.scala 31:69:@40077.4]
  wire [15:0] _T_95357; // @[Mux.scala 31:69:@40078.4]
  wire [15:0] _T_95358; // @[Mux.scala 31:69:@40079.4]
  wire [15:0] _T_95359; // @[Mux.scala 31:69:@40080.4]
  wire [15:0] _T_95360; // @[Mux.scala 31:69:@40081.4]
  wire [15:0] _T_95361; // @[Mux.scala 31:69:@40082.4]
  wire [15:0] _T_95362; // @[Mux.scala 31:69:@40083.4]
  wire [15:0] _T_95363; // @[Mux.scala 31:69:@40084.4]
  wire [15:0] _T_95364; // @[Mux.scala 31:69:@40085.4]
  wire [15:0] _T_95365; // @[Mux.scala 31:69:@40086.4]
  wire [15:0] _T_95366; // @[Mux.scala 31:69:@40087.4]
  wire [15:0] _T_95367; // @[Mux.scala 31:69:@40088.4]
  wire [15:0] _T_95368; // @[Mux.scala 31:69:@40089.4]
  wire [15:0] _T_95369; // @[Mux.scala 31:69:@40090.4]
  wire [15:0] _T_95370; // @[Mux.scala 31:69:@40091.4]
  wire [15:0] _T_95371; // @[Mux.scala 31:69:@40092.4]
  wire  _T_95372; // @[OneHot.scala 66:30:@40093.4]
  wire  _T_95373; // @[OneHot.scala 66:30:@40094.4]
  wire  _T_95374; // @[OneHot.scala 66:30:@40095.4]
  wire  _T_95375; // @[OneHot.scala 66:30:@40096.4]
  wire  _T_95376; // @[OneHot.scala 66:30:@40097.4]
  wire  _T_95377; // @[OneHot.scala 66:30:@40098.4]
  wire  _T_95378; // @[OneHot.scala 66:30:@40099.4]
  wire  _T_95379; // @[OneHot.scala 66:30:@40100.4]
  wire  _T_95380; // @[OneHot.scala 66:30:@40101.4]
  wire  _T_95381; // @[OneHot.scala 66:30:@40102.4]
  wire  _T_95382; // @[OneHot.scala 66:30:@40103.4]
  wire  _T_95383; // @[OneHot.scala 66:30:@40104.4]
  wire  _T_95384; // @[OneHot.scala 66:30:@40105.4]
  wire  _T_95385; // @[OneHot.scala 66:30:@40106.4]
  wire  _T_95386; // @[OneHot.scala 66:30:@40107.4]
  wire  _T_95387; // @[OneHot.scala 66:30:@40108.4]
  wire [15:0] _T_95428; // @[Mux.scala 31:69:@40126.4]
  wire [15:0] _T_95429; // @[Mux.scala 31:69:@40127.4]
  wire [15:0] _T_95430; // @[Mux.scala 31:69:@40128.4]
  wire [15:0] _T_95431; // @[Mux.scala 31:69:@40129.4]
  wire [15:0] _T_95432; // @[Mux.scala 31:69:@40130.4]
  wire [15:0] _T_95433; // @[Mux.scala 31:69:@40131.4]
  wire [15:0] _T_95434; // @[Mux.scala 31:69:@40132.4]
  wire [15:0] _T_95435; // @[Mux.scala 31:69:@40133.4]
  wire [15:0] _T_95436; // @[Mux.scala 31:69:@40134.4]
  wire [15:0] _T_95437; // @[Mux.scala 31:69:@40135.4]
  wire [15:0] _T_95438; // @[Mux.scala 31:69:@40136.4]
  wire [15:0] _T_95439; // @[Mux.scala 31:69:@40137.4]
  wire [15:0] _T_95440; // @[Mux.scala 31:69:@40138.4]
  wire [15:0] _T_95441; // @[Mux.scala 31:69:@40139.4]
  wire [15:0] _T_95442; // @[Mux.scala 31:69:@40140.4]
  wire [15:0] _T_95443; // @[Mux.scala 31:69:@40141.4]
  wire  _T_95444; // @[OneHot.scala 66:30:@40142.4]
  wire  _T_95445; // @[OneHot.scala 66:30:@40143.4]
  wire  _T_95446; // @[OneHot.scala 66:30:@40144.4]
  wire  _T_95447; // @[OneHot.scala 66:30:@40145.4]
  wire  _T_95448; // @[OneHot.scala 66:30:@40146.4]
  wire  _T_95449; // @[OneHot.scala 66:30:@40147.4]
  wire  _T_95450; // @[OneHot.scala 66:30:@40148.4]
  wire  _T_95451; // @[OneHot.scala 66:30:@40149.4]
  wire  _T_95452; // @[OneHot.scala 66:30:@40150.4]
  wire  _T_95453; // @[OneHot.scala 66:30:@40151.4]
  wire  _T_95454; // @[OneHot.scala 66:30:@40152.4]
  wire  _T_95455; // @[OneHot.scala 66:30:@40153.4]
  wire  _T_95456; // @[OneHot.scala 66:30:@40154.4]
  wire  _T_95457; // @[OneHot.scala 66:30:@40155.4]
  wire  _T_95458; // @[OneHot.scala 66:30:@40156.4]
  wire  _T_95459; // @[OneHot.scala 66:30:@40157.4]
  wire [15:0] _T_95500; // @[Mux.scala 31:69:@40175.4]
  wire [15:0] _T_95501; // @[Mux.scala 31:69:@40176.4]
  wire [15:0] _T_95502; // @[Mux.scala 31:69:@40177.4]
  wire [15:0] _T_95503; // @[Mux.scala 31:69:@40178.4]
  wire [15:0] _T_95504; // @[Mux.scala 31:69:@40179.4]
  wire [15:0] _T_95505; // @[Mux.scala 31:69:@40180.4]
  wire [15:0] _T_95506; // @[Mux.scala 31:69:@40181.4]
  wire [15:0] _T_95507; // @[Mux.scala 31:69:@40182.4]
  wire [15:0] _T_95508; // @[Mux.scala 31:69:@40183.4]
  wire [15:0] _T_95509; // @[Mux.scala 31:69:@40184.4]
  wire [15:0] _T_95510; // @[Mux.scala 31:69:@40185.4]
  wire [15:0] _T_95511; // @[Mux.scala 31:69:@40186.4]
  wire [15:0] _T_95512; // @[Mux.scala 31:69:@40187.4]
  wire [15:0] _T_95513; // @[Mux.scala 31:69:@40188.4]
  wire [15:0] _T_95514; // @[Mux.scala 31:69:@40189.4]
  wire [15:0] _T_95515; // @[Mux.scala 31:69:@40190.4]
  wire  _T_95516; // @[OneHot.scala 66:30:@40191.4]
  wire  _T_95517; // @[OneHot.scala 66:30:@40192.4]
  wire  _T_95518; // @[OneHot.scala 66:30:@40193.4]
  wire  _T_95519; // @[OneHot.scala 66:30:@40194.4]
  wire  _T_95520; // @[OneHot.scala 66:30:@40195.4]
  wire  _T_95521; // @[OneHot.scala 66:30:@40196.4]
  wire  _T_95522; // @[OneHot.scala 66:30:@40197.4]
  wire  _T_95523; // @[OneHot.scala 66:30:@40198.4]
  wire  _T_95524; // @[OneHot.scala 66:30:@40199.4]
  wire  _T_95525; // @[OneHot.scala 66:30:@40200.4]
  wire  _T_95526; // @[OneHot.scala 66:30:@40201.4]
  wire  _T_95527; // @[OneHot.scala 66:30:@40202.4]
  wire  _T_95528; // @[OneHot.scala 66:30:@40203.4]
  wire  _T_95529; // @[OneHot.scala 66:30:@40204.4]
  wire  _T_95530; // @[OneHot.scala 66:30:@40205.4]
  wire  _T_95531; // @[OneHot.scala 66:30:@40206.4]
  wire [15:0] _T_95572; // @[Mux.scala 31:69:@40224.4]
  wire [15:0] _T_95573; // @[Mux.scala 31:69:@40225.4]
  wire [15:0] _T_95574; // @[Mux.scala 31:69:@40226.4]
  wire [15:0] _T_95575; // @[Mux.scala 31:69:@40227.4]
  wire [15:0] _T_95576; // @[Mux.scala 31:69:@40228.4]
  wire [15:0] _T_95577; // @[Mux.scala 31:69:@40229.4]
  wire [15:0] _T_95578; // @[Mux.scala 31:69:@40230.4]
  wire [15:0] _T_95579; // @[Mux.scala 31:69:@40231.4]
  wire [15:0] _T_95580; // @[Mux.scala 31:69:@40232.4]
  wire [15:0] _T_95581; // @[Mux.scala 31:69:@40233.4]
  wire [15:0] _T_95582; // @[Mux.scala 31:69:@40234.4]
  wire [15:0] _T_95583; // @[Mux.scala 31:69:@40235.4]
  wire [15:0] _T_95584; // @[Mux.scala 31:69:@40236.4]
  wire [15:0] _T_95585; // @[Mux.scala 31:69:@40237.4]
  wire [15:0] _T_95586; // @[Mux.scala 31:69:@40238.4]
  wire [15:0] _T_95587; // @[Mux.scala 31:69:@40239.4]
  wire  _T_95588; // @[OneHot.scala 66:30:@40240.4]
  wire  _T_95589; // @[OneHot.scala 66:30:@40241.4]
  wire  _T_95590; // @[OneHot.scala 66:30:@40242.4]
  wire  _T_95591; // @[OneHot.scala 66:30:@40243.4]
  wire  _T_95592; // @[OneHot.scala 66:30:@40244.4]
  wire  _T_95593; // @[OneHot.scala 66:30:@40245.4]
  wire  _T_95594; // @[OneHot.scala 66:30:@40246.4]
  wire  _T_95595; // @[OneHot.scala 66:30:@40247.4]
  wire  _T_95596; // @[OneHot.scala 66:30:@40248.4]
  wire  _T_95597; // @[OneHot.scala 66:30:@40249.4]
  wire  _T_95598; // @[OneHot.scala 66:30:@40250.4]
  wire  _T_95599; // @[OneHot.scala 66:30:@40251.4]
  wire  _T_95600; // @[OneHot.scala 66:30:@40252.4]
  wire  _T_95601; // @[OneHot.scala 66:30:@40253.4]
  wire  _T_95602; // @[OneHot.scala 66:30:@40254.4]
  wire  _T_95603; // @[OneHot.scala 66:30:@40255.4]
  wire [15:0] _T_95644; // @[Mux.scala 31:69:@40273.4]
  wire [15:0] _T_95645; // @[Mux.scala 31:69:@40274.4]
  wire [15:0] _T_95646; // @[Mux.scala 31:69:@40275.4]
  wire [15:0] _T_95647; // @[Mux.scala 31:69:@40276.4]
  wire [15:0] _T_95648; // @[Mux.scala 31:69:@40277.4]
  wire [15:0] _T_95649; // @[Mux.scala 31:69:@40278.4]
  wire [15:0] _T_95650; // @[Mux.scala 31:69:@40279.4]
  wire [15:0] _T_95651; // @[Mux.scala 31:69:@40280.4]
  wire [15:0] _T_95652; // @[Mux.scala 31:69:@40281.4]
  wire [15:0] _T_95653; // @[Mux.scala 31:69:@40282.4]
  wire [15:0] _T_95654; // @[Mux.scala 31:69:@40283.4]
  wire [15:0] _T_95655; // @[Mux.scala 31:69:@40284.4]
  wire [15:0] _T_95656; // @[Mux.scala 31:69:@40285.4]
  wire [15:0] _T_95657; // @[Mux.scala 31:69:@40286.4]
  wire [15:0] _T_95658; // @[Mux.scala 31:69:@40287.4]
  wire [15:0] _T_95659; // @[Mux.scala 31:69:@40288.4]
  wire  _T_95660; // @[OneHot.scala 66:30:@40289.4]
  wire  _T_95661; // @[OneHot.scala 66:30:@40290.4]
  wire  _T_95662; // @[OneHot.scala 66:30:@40291.4]
  wire  _T_95663; // @[OneHot.scala 66:30:@40292.4]
  wire  _T_95664; // @[OneHot.scala 66:30:@40293.4]
  wire  _T_95665; // @[OneHot.scala 66:30:@40294.4]
  wire  _T_95666; // @[OneHot.scala 66:30:@40295.4]
  wire  _T_95667; // @[OneHot.scala 66:30:@40296.4]
  wire  _T_95668; // @[OneHot.scala 66:30:@40297.4]
  wire  _T_95669; // @[OneHot.scala 66:30:@40298.4]
  wire  _T_95670; // @[OneHot.scala 66:30:@40299.4]
  wire  _T_95671; // @[OneHot.scala 66:30:@40300.4]
  wire  _T_95672; // @[OneHot.scala 66:30:@40301.4]
  wire  _T_95673; // @[OneHot.scala 66:30:@40302.4]
  wire  _T_95674; // @[OneHot.scala 66:30:@40303.4]
  wire  _T_95675; // @[OneHot.scala 66:30:@40304.4]
  wire [7:0] _T_95740; // @[Mux.scala 19:72:@40328.4]
  wire [15:0] _T_95748; // @[Mux.scala 19:72:@40336.4]
  wire [15:0] _T_95750; // @[Mux.scala 19:72:@40337.4]
  wire [7:0] _T_95757; // @[Mux.scala 19:72:@40344.4]
  wire [15:0] _T_95765; // @[Mux.scala 19:72:@40352.4]
  wire [15:0] _T_95767; // @[Mux.scala 19:72:@40353.4]
  wire [7:0] _T_95774; // @[Mux.scala 19:72:@40360.4]
  wire [15:0] _T_95782; // @[Mux.scala 19:72:@40368.4]
  wire [15:0] _T_95784; // @[Mux.scala 19:72:@40369.4]
  wire [7:0] _T_95791; // @[Mux.scala 19:72:@40376.4]
  wire [15:0] _T_95799; // @[Mux.scala 19:72:@40384.4]
  wire [15:0] _T_95801; // @[Mux.scala 19:72:@40385.4]
  wire [7:0] _T_95808; // @[Mux.scala 19:72:@40392.4]
  wire [15:0] _T_95816; // @[Mux.scala 19:72:@40400.4]
  wire [15:0] _T_95818; // @[Mux.scala 19:72:@40401.4]
  wire [7:0] _T_95825; // @[Mux.scala 19:72:@40408.4]
  wire [15:0] _T_95833; // @[Mux.scala 19:72:@40416.4]
  wire [15:0] _T_95835; // @[Mux.scala 19:72:@40417.4]
  wire [7:0] _T_95842; // @[Mux.scala 19:72:@40424.4]
  wire [15:0] _T_95850; // @[Mux.scala 19:72:@40432.4]
  wire [15:0] _T_95852; // @[Mux.scala 19:72:@40433.4]
  wire [7:0] _T_95859; // @[Mux.scala 19:72:@40440.4]
  wire [15:0] _T_95867; // @[Mux.scala 19:72:@40448.4]
  wire [15:0] _T_95869; // @[Mux.scala 19:72:@40449.4]
  wire [7:0] _T_95876; // @[Mux.scala 19:72:@40456.4]
  wire [15:0] _T_95884; // @[Mux.scala 19:72:@40464.4]
  wire [15:0] _T_95886; // @[Mux.scala 19:72:@40465.4]
  wire [7:0] _T_95893; // @[Mux.scala 19:72:@40472.4]
  wire [15:0] _T_95901; // @[Mux.scala 19:72:@40480.4]
  wire [15:0] _T_95903; // @[Mux.scala 19:72:@40481.4]
  wire [7:0] _T_95910; // @[Mux.scala 19:72:@40488.4]
  wire [15:0] _T_95918; // @[Mux.scala 19:72:@40496.4]
  wire [15:0] _T_95920; // @[Mux.scala 19:72:@40497.4]
  wire [7:0] _T_95927; // @[Mux.scala 19:72:@40504.4]
  wire [15:0] _T_95935; // @[Mux.scala 19:72:@40512.4]
  wire [15:0] _T_95937; // @[Mux.scala 19:72:@40513.4]
  wire [7:0] _T_95944; // @[Mux.scala 19:72:@40520.4]
  wire [15:0] _T_95952; // @[Mux.scala 19:72:@40528.4]
  wire [15:0] _T_95954; // @[Mux.scala 19:72:@40529.4]
  wire [7:0] _T_95961; // @[Mux.scala 19:72:@40536.4]
  wire [15:0] _T_95969; // @[Mux.scala 19:72:@40544.4]
  wire [15:0] _T_95971; // @[Mux.scala 19:72:@40545.4]
  wire [7:0] _T_95978; // @[Mux.scala 19:72:@40552.4]
  wire [15:0] _T_95986; // @[Mux.scala 19:72:@40560.4]
  wire [15:0] _T_95988; // @[Mux.scala 19:72:@40561.4]
  wire [7:0] _T_95995; // @[Mux.scala 19:72:@40568.4]
  wire [15:0] _T_96003; // @[Mux.scala 19:72:@40576.4]
  wire [15:0] _T_96005; // @[Mux.scala 19:72:@40577.4]
  wire [15:0] _T_96006; // @[Mux.scala 19:72:@40578.4]
  wire [15:0] _T_96007; // @[Mux.scala 19:72:@40579.4]
  wire [15:0] _T_96008; // @[Mux.scala 19:72:@40580.4]
  wire [15:0] _T_96009; // @[Mux.scala 19:72:@40581.4]
  wire [15:0] _T_96010; // @[Mux.scala 19:72:@40582.4]
  wire [15:0] _T_96011; // @[Mux.scala 19:72:@40583.4]
  wire [15:0] _T_96012; // @[Mux.scala 19:72:@40584.4]
  wire [15:0] _T_96013; // @[Mux.scala 19:72:@40585.4]
  wire [15:0] _T_96014; // @[Mux.scala 19:72:@40586.4]
  wire [15:0] _T_96015; // @[Mux.scala 19:72:@40587.4]
  wire [15:0] _T_96016; // @[Mux.scala 19:72:@40588.4]
  wire [15:0] _T_96017; // @[Mux.scala 19:72:@40589.4]
  wire [15:0] _T_96018; // @[Mux.scala 19:72:@40590.4]
  wire [15:0] _T_96019; // @[Mux.scala 19:72:@40591.4]
  wire [15:0] _T_96020; // @[Mux.scala 19:72:@40592.4]
  wire  inputPriorityPorts_0_0; // @[Mux.scala 19:72:@40596.4]
  wire  inputPriorityPorts_0_1; // @[Mux.scala 19:72:@40598.4]
  wire  inputPriorityPorts_0_2; // @[Mux.scala 19:72:@40600.4]
  wire  inputPriorityPorts_0_3; // @[Mux.scala 19:72:@40602.4]
  wire  inputPriorityPorts_0_4; // @[Mux.scala 19:72:@40604.4]
  wire  inputPriorityPorts_0_5; // @[Mux.scala 19:72:@40606.4]
  wire  inputPriorityPorts_0_6; // @[Mux.scala 19:72:@40608.4]
  wire  inputPriorityPorts_0_7; // @[Mux.scala 19:72:@40610.4]
  wire  inputPriorityPorts_0_8; // @[Mux.scala 19:72:@40612.4]
  wire  inputPriorityPorts_0_9; // @[Mux.scala 19:72:@40614.4]
  wire  inputPriorityPorts_0_10; // @[Mux.scala 19:72:@40616.4]
  wire  inputPriorityPorts_0_11; // @[Mux.scala 19:72:@40618.4]
  wire  inputPriorityPorts_0_12; // @[Mux.scala 19:72:@40620.4]
  wire  inputPriorityPorts_0_13; // @[Mux.scala 19:72:@40622.4]
  wire  inputPriorityPorts_0_14; // @[Mux.scala 19:72:@40624.4]
  wire  inputPriorityPorts_0_15; // @[Mux.scala 19:72:@40626.4]
  wire [15:0] _T_96222; // @[Mux.scala 31:69:@40680.4]
  wire [15:0] _T_96223; // @[Mux.scala 31:69:@40681.4]
  wire [15:0] _T_96224; // @[Mux.scala 31:69:@40682.4]
  wire [15:0] _T_96225; // @[Mux.scala 31:69:@40683.4]
  wire [15:0] _T_96226; // @[Mux.scala 31:69:@40684.4]
  wire [15:0] _T_96227; // @[Mux.scala 31:69:@40685.4]
  wire [15:0] _T_96228; // @[Mux.scala 31:69:@40686.4]
  wire [15:0] _T_96229; // @[Mux.scala 31:69:@40687.4]
  wire [15:0] _T_96230; // @[Mux.scala 31:69:@40688.4]
  wire [15:0] _T_96231; // @[Mux.scala 31:69:@40689.4]
  wire [15:0] _T_96232; // @[Mux.scala 31:69:@40690.4]
  wire [15:0] _T_96233; // @[Mux.scala 31:69:@40691.4]
  wire [15:0] _T_96234; // @[Mux.scala 31:69:@40692.4]
  wire [15:0] _T_96235; // @[Mux.scala 31:69:@40693.4]
  wire [15:0] _T_96236; // @[Mux.scala 31:69:@40694.4]
  wire [15:0] _T_96237; // @[Mux.scala 31:69:@40695.4]
  wire  _T_96238; // @[OneHot.scala 66:30:@40696.4]
  wire  _T_96239; // @[OneHot.scala 66:30:@40697.4]
  wire  _T_96240; // @[OneHot.scala 66:30:@40698.4]
  wire  _T_96241; // @[OneHot.scala 66:30:@40699.4]
  wire  _T_96242; // @[OneHot.scala 66:30:@40700.4]
  wire  _T_96243; // @[OneHot.scala 66:30:@40701.4]
  wire  _T_96244; // @[OneHot.scala 66:30:@40702.4]
  wire  _T_96245; // @[OneHot.scala 66:30:@40703.4]
  wire  _T_96246; // @[OneHot.scala 66:30:@40704.4]
  wire  _T_96247; // @[OneHot.scala 66:30:@40705.4]
  wire  _T_96248; // @[OneHot.scala 66:30:@40706.4]
  wire  _T_96249; // @[OneHot.scala 66:30:@40707.4]
  wire  _T_96250; // @[OneHot.scala 66:30:@40708.4]
  wire  _T_96251; // @[OneHot.scala 66:30:@40709.4]
  wire  _T_96252; // @[OneHot.scala 66:30:@40710.4]
  wire  _T_96253; // @[OneHot.scala 66:30:@40711.4]
  wire [15:0] _T_96294; // @[Mux.scala 31:69:@40729.4]
  wire [15:0] _T_96295; // @[Mux.scala 31:69:@40730.4]
  wire [15:0] _T_96296; // @[Mux.scala 31:69:@40731.4]
  wire [15:0] _T_96297; // @[Mux.scala 31:69:@40732.4]
  wire [15:0] _T_96298; // @[Mux.scala 31:69:@40733.4]
  wire [15:0] _T_96299; // @[Mux.scala 31:69:@40734.4]
  wire [15:0] _T_96300; // @[Mux.scala 31:69:@40735.4]
  wire [15:0] _T_96301; // @[Mux.scala 31:69:@40736.4]
  wire [15:0] _T_96302; // @[Mux.scala 31:69:@40737.4]
  wire [15:0] _T_96303; // @[Mux.scala 31:69:@40738.4]
  wire [15:0] _T_96304; // @[Mux.scala 31:69:@40739.4]
  wire [15:0] _T_96305; // @[Mux.scala 31:69:@40740.4]
  wire [15:0] _T_96306; // @[Mux.scala 31:69:@40741.4]
  wire [15:0] _T_96307; // @[Mux.scala 31:69:@40742.4]
  wire [15:0] _T_96308; // @[Mux.scala 31:69:@40743.4]
  wire [15:0] _T_96309; // @[Mux.scala 31:69:@40744.4]
  wire  _T_96310; // @[OneHot.scala 66:30:@40745.4]
  wire  _T_96311; // @[OneHot.scala 66:30:@40746.4]
  wire  _T_96312; // @[OneHot.scala 66:30:@40747.4]
  wire  _T_96313; // @[OneHot.scala 66:30:@40748.4]
  wire  _T_96314; // @[OneHot.scala 66:30:@40749.4]
  wire  _T_96315; // @[OneHot.scala 66:30:@40750.4]
  wire  _T_96316; // @[OneHot.scala 66:30:@40751.4]
  wire  _T_96317; // @[OneHot.scala 66:30:@40752.4]
  wire  _T_96318; // @[OneHot.scala 66:30:@40753.4]
  wire  _T_96319; // @[OneHot.scala 66:30:@40754.4]
  wire  _T_96320; // @[OneHot.scala 66:30:@40755.4]
  wire  _T_96321; // @[OneHot.scala 66:30:@40756.4]
  wire  _T_96322; // @[OneHot.scala 66:30:@40757.4]
  wire  _T_96323; // @[OneHot.scala 66:30:@40758.4]
  wire  _T_96324; // @[OneHot.scala 66:30:@40759.4]
  wire  _T_96325; // @[OneHot.scala 66:30:@40760.4]
  wire [15:0] _T_96366; // @[Mux.scala 31:69:@40778.4]
  wire [15:0] _T_96367; // @[Mux.scala 31:69:@40779.4]
  wire [15:0] _T_96368; // @[Mux.scala 31:69:@40780.4]
  wire [15:0] _T_96369; // @[Mux.scala 31:69:@40781.4]
  wire [15:0] _T_96370; // @[Mux.scala 31:69:@40782.4]
  wire [15:0] _T_96371; // @[Mux.scala 31:69:@40783.4]
  wire [15:0] _T_96372; // @[Mux.scala 31:69:@40784.4]
  wire [15:0] _T_96373; // @[Mux.scala 31:69:@40785.4]
  wire [15:0] _T_96374; // @[Mux.scala 31:69:@40786.4]
  wire [15:0] _T_96375; // @[Mux.scala 31:69:@40787.4]
  wire [15:0] _T_96376; // @[Mux.scala 31:69:@40788.4]
  wire [15:0] _T_96377; // @[Mux.scala 31:69:@40789.4]
  wire [15:0] _T_96378; // @[Mux.scala 31:69:@40790.4]
  wire [15:0] _T_96379; // @[Mux.scala 31:69:@40791.4]
  wire [15:0] _T_96380; // @[Mux.scala 31:69:@40792.4]
  wire [15:0] _T_96381; // @[Mux.scala 31:69:@40793.4]
  wire  _T_96382; // @[OneHot.scala 66:30:@40794.4]
  wire  _T_96383; // @[OneHot.scala 66:30:@40795.4]
  wire  _T_96384; // @[OneHot.scala 66:30:@40796.4]
  wire  _T_96385; // @[OneHot.scala 66:30:@40797.4]
  wire  _T_96386; // @[OneHot.scala 66:30:@40798.4]
  wire  _T_96387; // @[OneHot.scala 66:30:@40799.4]
  wire  _T_96388; // @[OneHot.scala 66:30:@40800.4]
  wire  _T_96389; // @[OneHot.scala 66:30:@40801.4]
  wire  _T_96390; // @[OneHot.scala 66:30:@40802.4]
  wire  _T_96391; // @[OneHot.scala 66:30:@40803.4]
  wire  _T_96392; // @[OneHot.scala 66:30:@40804.4]
  wire  _T_96393; // @[OneHot.scala 66:30:@40805.4]
  wire  _T_96394; // @[OneHot.scala 66:30:@40806.4]
  wire  _T_96395; // @[OneHot.scala 66:30:@40807.4]
  wire  _T_96396; // @[OneHot.scala 66:30:@40808.4]
  wire  _T_96397; // @[OneHot.scala 66:30:@40809.4]
  wire [15:0] _T_96438; // @[Mux.scala 31:69:@40827.4]
  wire [15:0] _T_96439; // @[Mux.scala 31:69:@40828.4]
  wire [15:0] _T_96440; // @[Mux.scala 31:69:@40829.4]
  wire [15:0] _T_96441; // @[Mux.scala 31:69:@40830.4]
  wire [15:0] _T_96442; // @[Mux.scala 31:69:@40831.4]
  wire [15:0] _T_96443; // @[Mux.scala 31:69:@40832.4]
  wire [15:0] _T_96444; // @[Mux.scala 31:69:@40833.4]
  wire [15:0] _T_96445; // @[Mux.scala 31:69:@40834.4]
  wire [15:0] _T_96446; // @[Mux.scala 31:69:@40835.4]
  wire [15:0] _T_96447; // @[Mux.scala 31:69:@40836.4]
  wire [15:0] _T_96448; // @[Mux.scala 31:69:@40837.4]
  wire [15:0] _T_96449; // @[Mux.scala 31:69:@40838.4]
  wire [15:0] _T_96450; // @[Mux.scala 31:69:@40839.4]
  wire [15:0] _T_96451; // @[Mux.scala 31:69:@40840.4]
  wire [15:0] _T_96452; // @[Mux.scala 31:69:@40841.4]
  wire [15:0] _T_96453; // @[Mux.scala 31:69:@40842.4]
  wire  _T_96454; // @[OneHot.scala 66:30:@40843.4]
  wire  _T_96455; // @[OneHot.scala 66:30:@40844.4]
  wire  _T_96456; // @[OneHot.scala 66:30:@40845.4]
  wire  _T_96457; // @[OneHot.scala 66:30:@40846.4]
  wire  _T_96458; // @[OneHot.scala 66:30:@40847.4]
  wire  _T_96459; // @[OneHot.scala 66:30:@40848.4]
  wire  _T_96460; // @[OneHot.scala 66:30:@40849.4]
  wire  _T_96461; // @[OneHot.scala 66:30:@40850.4]
  wire  _T_96462; // @[OneHot.scala 66:30:@40851.4]
  wire  _T_96463; // @[OneHot.scala 66:30:@40852.4]
  wire  _T_96464; // @[OneHot.scala 66:30:@40853.4]
  wire  _T_96465; // @[OneHot.scala 66:30:@40854.4]
  wire  _T_96466; // @[OneHot.scala 66:30:@40855.4]
  wire  _T_96467; // @[OneHot.scala 66:30:@40856.4]
  wire  _T_96468; // @[OneHot.scala 66:30:@40857.4]
  wire  _T_96469; // @[OneHot.scala 66:30:@40858.4]
  wire [15:0] _T_96510; // @[Mux.scala 31:69:@40876.4]
  wire [15:0] _T_96511; // @[Mux.scala 31:69:@40877.4]
  wire [15:0] _T_96512; // @[Mux.scala 31:69:@40878.4]
  wire [15:0] _T_96513; // @[Mux.scala 31:69:@40879.4]
  wire [15:0] _T_96514; // @[Mux.scala 31:69:@40880.4]
  wire [15:0] _T_96515; // @[Mux.scala 31:69:@40881.4]
  wire [15:0] _T_96516; // @[Mux.scala 31:69:@40882.4]
  wire [15:0] _T_96517; // @[Mux.scala 31:69:@40883.4]
  wire [15:0] _T_96518; // @[Mux.scala 31:69:@40884.4]
  wire [15:0] _T_96519; // @[Mux.scala 31:69:@40885.4]
  wire [15:0] _T_96520; // @[Mux.scala 31:69:@40886.4]
  wire [15:0] _T_96521; // @[Mux.scala 31:69:@40887.4]
  wire [15:0] _T_96522; // @[Mux.scala 31:69:@40888.4]
  wire [15:0] _T_96523; // @[Mux.scala 31:69:@40889.4]
  wire [15:0] _T_96524; // @[Mux.scala 31:69:@40890.4]
  wire [15:0] _T_96525; // @[Mux.scala 31:69:@40891.4]
  wire  _T_96526; // @[OneHot.scala 66:30:@40892.4]
  wire  _T_96527; // @[OneHot.scala 66:30:@40893.4]
  wire  _T_96528; // @[OneHot.scala 66:30:@40894.4]
  wire  _T_96529; // @[OneHot.scala 66:30:@40895.4]
  wire  _T_96530; // @[OneHot.scala 66:30:@40896.4]
  wire  _T_96531; // @[OneHot.scala 66:30:@40897.4]
  wire  _T_96532; // @[OneHot.scala 66:30:@40898.4]
  wire  _T_96533; // @[OneHot.scala 66:30:@40899.4]
  wire  _T_96534; // @[OneHot.scala 66:30:@40900.4]
  wire  _T_96535; // @[OneHot.scala 66:30:@40901.4]
  wire  _T_96536; // @[OneHot.scala 66:30:@40902.4]
  wire  _T_96537; // @[OneHot.scala 66:30:@40903.4]
  wire  _T_96538; // @[OneHot.scala 66:30:@40904.4]
  wire  _T_96539; // @[OneHot.scala 66:30:@40905.4]
  wire  _T_96540; // @[OneHot.scala 66:30:@40906.4]
  wire  _T_96541; // @[OneHot.scala 66:30:@40907.4]
  wire [15:0] _T_96582; // @[Mux.scala 31:69:@40925.4]
  wire [15:0] _T_96583; // @[Mux.scala 31:69:@40926.4]
  wire [15:0] _T_96584; // @[Mux.scala 31:69:@40927.4]
  wire [15:0] _T_96585; // @[Mux.scala 31:69:@40928.4]
  wire [15:0] _T_96586; // @[Mux.scala 31:69:@40929.4]
  wire [15:0] _T_96587; // @[Mux.scala 31:69:@40930.4]
  wire [15:0] _T_96588; // @[Mux.scala 31:69:@40931.4]
  wire [15:0] _T_96589; // @[Mux.scala 31:69:@40932.4]
  wire [15:0] _T_96590; // @[Mux.scala 31:69:@40933.4]
  wire [15:0] _T_96591; // @[Mux.scala 31:69:@40934.4]
  wire [15:0] _T_96592; // @[Mux.scala 31:69:@40935.4]
  wire [15:0] _T_96593; // @[Mux.scala 31:69:@40936.4]
  wire [15:0] _T_96594; // @[Mux.scala 31:69:@40937.4]
  wire [15:0] _T_96595; // @[Mux.scala 31:69:@40938.4]
  wire [15:0] _T_96596; // @[Mux.scala 31:69:@40939.4]
  wire [15:0] _T_96597; // @[Mux.scala 31:69:@40940.4]
  wire  _T_96598; // @[OneHot.scala 66:30:@40941.4]
  wire  _T_96599; // @[OneHot.scala 66:30:@40942.4]
  wire  _T_96600; // @[OneHot.scala 66:30:@40943.4]
  wire  _T_96601; // @[OneHot.scala 66:30:@40944.4]
  wire  _T_96602; // @[OneHot.scala 66:30:@40945.4]
  wire  _T_96603; // @[OneHot.scala 66:30:@40946.4]
  wire  _T_96604; // @[OneHot.scala 66:30:@40947.4]
  wire  _T_96605; // @[OneHot.scala 66:30:@40948.4]
  wire  _T_96606; // @[OneHot.scala 66:30:@40949.4]
  wire  _T_96607; // @[OneHot.scala 66:30:@40950.4]
  wire  _T_96608; // @[OneHot.scala 66:30:@40951.4]
  wire  _T_96609; // @[OneHot.scala 66:30:@40952.4]
  wire  _T_96610; // @[OneHot.scala 66:30:@40953.4]
  wire  _T_96611; // @[OneHot.scala 66:30:@40954.4]
  wire  _T_96612; // @[OneHot.scala 66:30:@40955.4]
  wire  _T_96613; // @[OneHot.scala 66:30:@40956.4]
  wire [15:0] _T_96654; // @[Mux.scala 31:69:@40974.4]
  wire [15:0] _T_96655; // @[Mux.scala 31:69:@40975.4]
  wire [15:0] _T_96656; // @[Mux.scala 31:69:@40976.4]
  wire [15:0] _T_96657; // @[Mux.scala 31:69:@40977.4]
  wire [15:0] _T_96658; // @[Mux.scala 31:69:@40978.4]
  wire [15:0] _T_96659; // @[Mux.scala 31:69:@40979.4]
  wire [15:0] _T_96660; // @[Mux.scala 31:69:@40980.4]
  wire [15:0] _T_96661; // @[Mux.scala 31:69:@40981.4]
  wire [15:0] _T_96662; // @[Mux.scala 31:69:@40982.4]
  wire [15:0] _T_96663; // @[Mux.scala 31:69:@40983.4]
  wire [15:0] _T_96664; // @[Mux.scala 31:69:@40984.4]
  wire [15:0] _T_96665; // @[Mux.scala 31:69:@40985.4]
  wire [15:0] _T_96666; // @[Mux.scala 31:69:@40986.4]
  wire [15:0] _T_96667; // @[Mux.scala 31:69:@40987.4]
  wire [15:0] _T_96668; // @[Mux.scala 31:69:@40988.4]
  wire [15:0] _T_96669; // @[Mux.scala 31:69:@40989.4]
  wire  _T_96670; // @[OneHot.scala 66:30:@40990.4]
  wire  _T_96671; // @[OneHot.scala 66:30:@40991.4]
  wire  _T_96672; // @[OneHot.scala 66:30:@40992.4]
  wire  _T_96673; // @[OneHot.scala 66:30:@40993.4]
  wire  _T_96674; // @[OneHot.scala 66:30:@40994.4]
  wire  _T_96675; // @[OneHot.scala 66:30:@40995.4]
  wire  _T_96676; // @[OneHot.scala 66:30:@40996.4]
  wire  _T_96677; // @[OneHot.scala 66:30:@40997.4]
  wire  _T_96678; // @[OneHot.scala 66:30:@40998.4]
  wire  _T_96679; // @[OneHot.scala 66:30:@40999.4]
  wire  _T_96680; // @[OneHot.scala 66:30:@41000.4]
  wire  _T_96681; // @[OneHot.scala 66:30:@41001.4]
  wire  _T_96682; // @[OneHot.scala 66:30:@41002.4]
  wire  _T_96683; // @[OneHot.scala 66:30:@41003.4]
  wire  _T_96684; // @[OneHot.scala 66:30:@41004.4]
  wire  _T_96685; // @[OneHot.scala 66:30:@41005.4]
  wire [15:0] _T_96726; // @[Mux.scala 31:69:@41023.4]
  wire [15:0] _T_96727; // @[Mux.scala 31:69:@41024.4]
  wire [15:0] _T_96728; // @[Mux.scala 31:69:@41025.4]
  wire [15:0] _T_96729; // @[Mux.scala 31:69:@41026.4]
  wire [15:0] _T_96730; // @[Mux.scala 31:69:@41027.4]
  wire [15:0] _T_96731; // @[Mux.scala 31:69:@41028.4]
  wire [15:0] _T_96732; // @[Mux.scala 31:69:@41029.4]
  wire [15:0] _T_96733; // @[Mux.scala 31:69:@41030.4]
  wire [15:0] _T_96734; // @[Mux.scala 31:69:@41031.4]
  wire [15:0] _T_96735; // @[Mux.scala 31:69:@41032.4]
  wire [15:0] _T_96736; // @[Mux.scala 31:69:@41033.4]
  wire [15:0] _T_96737; // @[Mux.scala 31:69:@41034.4]
  wire [15:0] _T_96738; // @[Mux.scala 31:69:@41035.4]
  wire [15:0] _T_96739; // @[Mux.scala 31:69:@41036.4]
  wire [15:0] _T_96740; // @[Mux.scala 31:69:@41037.4]
  wire [15:0] _T_96741; // @[Mux.scala 31:69:@41038.4]
  wire  _T_96742; // @[OneHot.scala 66:30:@41039.4]
  wire  _T_96743; // @[OneHot.scala 66:30:@41040.4]
  wire  _T_96744; // @[OneHot.scala 66:30:@41041.4]
  wire  _T_96745; // @[OneHot.scala 66:30:@41042.4]
  wire  _T_96746; // @[OneHot.scala 66:30:@41043.4]
  wire  _T_96747; // @[OneHot.scala 66:30:@41044.4]
  wire  _T_96748; // @[OneHot.scala 66:30:@41045.4]
  wire  _T_96749; // @[OneHot.scala 66:30:@41046.4]
  wire  _T_96750; // @[OneHot.scala 66:30:@41047.4]
  wire  _T_96751; // @[OneHot.scala 66:30:@41048.4]
  wire  _T_96752; // @[OneHot.scala 66:30:@41049.4]
  wire  _T_96753; // @[OneHot.scala 66:30:@41050.4]
  wire  _T_96754; // @[OneHot.scala 66:30:@41051.4]
  wire  _T_96755; // @[OneHot.scala 66:30:@41052.4]
  wire  _T_96756; // @[OneHot.scala 66:30:@41053.4]
  wire  _T_96757; // @[OneHot.scala 66:30:@41054.4]
  wire [15:0] _T_96798; // @[Mux.scala 31:69:@41072.4]
  wire [15:0] _T_96799; // @[Mux.scala 31:69:@41073.4]
  wire [15:0] _T_96800; // @[Mux.scala 31:69:@41074.4]
  wire [15:0] _T_96801; // @[Mux.scala 31:69:@41075.4]
  wire [15:0] _T_96802; // @[Mux.scala 31:69:@41076.4]
  wire [15:0] _T_96803; // @[Mux.scala 31:69:@41077.4]
  wire [15:0] _T_96804; // @[Mux.scala 31:69:@41078.4]
  wire [15:0] _T_96805; // @[Mux.scala 31:69:@41079.4]
  wire [15:0] _T_96806; // @[Mux.scala 31:69:@41080.4]
  wire [15:0] _T_96807; // @[Mux.scala 31:69:@41081.4]
  wire [15:0] _T_96808; // @[Mux.scala 31:69:@41082.4]
  wire [15:0] _T_96809; // @[Mux.scala 31:69:@41083.4]
  wire [15:0] _T_96810; // @[Mux.scala 31:69:@41084.4]
  wire [15:0] _T_96811; // @[Mux.scala 31:69:@41085.4]
  wire [15:0] _T_96812; // @[Mux.scala 31:69:@41086.4]
  wire [15:0] _T_96813; // @[Mux.scala 31:69:@41087.4]
  wire  _T_96814; // @[OneHot.scala 66:30:@41088.4]
  wire  _T_96815; // @[OneHot.scala 66:30:@41089.4]
  wire  _T_96816; // @[OneHot.scala 66:30:@41090.4]
  wire  _T_96817; // @[OneHot.scala 66:30:@41091.4]
  wire  _T_96818; // @[OneHot.scala 66:30:@41092.4]
  wire  _T_96819; // @[OneHot.scala 66:30:@41093.4]
  wire  _T_96820; // @[OneHot.scala 66:30:@41094.4]
  wire  _T_96821; // @[OneHot.scala 66:30:@41095.4]
  wire  _T_96822; // @[OneHot.scala 66:30:@41096.4]
  wire  _T_96823; // @[OneHot.scala 66:30:@41097.4]
  wire  _T_96824; // @[OneHot.scala 66:30:@41098.4]
  wire  _T_96825; // @[OneHot.scala 66:30:@41099.4]
  wire  _T_96826; // @[OneHot.scala 66:30:@41100.4]
  wire  _T_96827; // @[OneHot.scala 66:30:@41101.4]
  wire  _T_96828; // @[OneHot.scala 66:30:@41102.4]
  wire  _T_96829; // @[OneHot.scala 66:30:@41103.4]
  wire [15:0] _T_96870; // @[Mux.scala 31:69:@41121.4]
  wire [15:0] _T_96871; // @[Mux.scala 31:69:@41122.4]
  wire [15:0] _T_96872; // @[Mux.scala 31:69:@41123.4]
  wire [15:0] _T_96873; // @[Mux.scala 31:69:@41124.4]
  wire [15:0] _T_96874; // @[Mux.scala 31:69:@41125.4]
  wire [15:0] _T_96875; // @[Mux.scala 31:69:@41126.4]
  wire [15:0] _T_96876; // @[Mux.scala 31:69:@41127.4]
  wire [15:0] _T_96877; // @[Mux.scala 31:69:@41128.4]
  wire [15:0] _T_96878; // @[Mux.scala 31:69:@41129.4]
  wire [15:0] _T_96879; // @[Mux.scala 31:69:@41130.4]
  wire [15:0] _T_96880; // @[Mux.scala 31:69:@41131.4]
  wire [15:0] _T_96881; // @[Mux.scala 31:69:@41132.4]
  wire [15:0] _T_96882; // @[Mux.scala 31:69:@41133.4]
  wire [15:0] _T_96883; // @[Mux.scala 31:69:@41134.4]
  wire [15:0] _T_96884; // @[Mux.scala 31:69:@41135.4]
  wire [15:0] _T_96885; // @[Mux.scala 31:69:@41136.4]
  wire  _T_96886; // @[OneHot.scala 66:30:@41137.4]
  wire  _T_96887; // @[OneHot.scala 66:30:@41138.4]
  wire  _T_96888; // @[OneHot.scala 66:30:@41139.4]
  wire  _T_96889; // @[OneHot.scala 66:30:@41140.4]
  wire  _T_96890; // @[OneHot.scala 66:30:@41141.4]
  wire  _T_96891; // @[OneHot.scala 66:30:@41142.4]
  wire  _T_96892; // @[OneHot.scala 66:30:@41143.4]
  wire  _T_96893; // @[OneHot.scala 66:30:@41144.4]
  wire  _T_96894; // @[OneHot.scala 66:30:@41145.4]
  wire  _T_96895; // @[OneHot.scala 66:30:@41146.4]
  wire  _T_96896; // @[OneHot.scala 66:30:@41147.4]
  wire  _T_96897; // @[OneHot.scala 66:30:@41148.4]
  wire  _T_96898; // @[OneHot.scala 66:30:@41149.4]
  wire  _T_96899; // @[OneHot.scala 66:30:@41150.4]
  wire  _T_96900; // @[OneHot.scala 66:30:@41151.4]
  wire  _T_96901; // @[OneHot.scala 66:30:@41152.4]
  wire [15:0] _T_96942; // @[Mux.scala 31:69:@41170.4]
  wire [15:0] _T_96943; // @[Mux.scala 31:69:@41171.4]
  wire [15:0] _T_96944; // @[Mux.scala 31:69:@41172.4]
  wire [15:0] _T_96945; // @[Mux.scala 31:69:@41173.4]
  wire [15:0] _T_96946; // @[Mux.scala 31:69:@41174.4]
  wire [15:0] _T_96947; // @[Mux.scala 31:69:@41175.4]
  wire [15:0] _T_96948; // @[Mux.scala 31:69:@41176.4]
  wire [15:0] _T_96949; // @[Mux.scala 31:69:@41177.4]
  wire [15:0] _T_96950; // @[Mux.scala 31:69:@41178.4]
  wire [15:0] _T_96951; // @[Mux.scala 31:69:@41179.4]
  wire [15:0] _T_96952; // @[Mux.scala 31:69:@41180.4]
  wire [15:0] _T_96953; // @[Mux.scala 31:69:@41181.4]
  wire [15:0] _T_96954; // @[Mux.scala 31:69:@41182.4]
  wire [15:0] _T_96955; // @[Mux.scala 31:69:@41183.4]
  wire [15:0] _T_96956; // @[Mux.scala 31:69:@41184.4]
  wire [15:0] _T_96957; // @[Mux.scala 31:69:@41185.4]
  wire  _T_96958; // @[OneHot.scala 66:30:@41186.4]
  wire  _T_96959; // @[OneHot.scala 66:30:@41187.4]
  wire  _T_96960; // @[OneHot.scala 66:30:@41188.4]
  wire  _T_96961; // @[OneHot.scala 66:30:@41189.4]
  wire  _T_96962; // @[OneHot.scala 66:30:@41190.4]
  wire  _T_96963; // @[OneHot.scala 66:30:@41191.4]
  wire  _T_96964; // @[OneHot.scala 66:30:@41192.4]
  wire  _T_96965; // @[OneHot.scala 66:30:@41193.4]
  wire  _T_96966; // @[OneHot.scala 66:30:@41194.4]
  wire  _T_96967; // @[OneHot.scala 66:30:@41195.4]
  wire  _T_96968; // @[OneHot.scala 66:30:@41196.4]
  wire  _T_96969; // @[OneHot.scala 66:30:@41197.4]
  wire  _T_96970; // @[OneHot.scala 66:30:@41198.4]
  wire  _T_96971; // @[OneHot.scala 66:30:@41199.4]
  wire  _T_96972; // @[OneHot.scala 66:30:@41200.4]
  wire  _T_96973; // @[OneHot.scala 66:30:@41201.4]
  wire [15:0] _T_97014; // @[Mux.scala 31:69:@41219.4]
  wire [15:0] _T_97015; // @[Mux.scala 31:69:@41220.4]
  wire [15:0] _T_97016; // @[Mux.scala 31:69:@41221.4]
  wire [15:0] _T_97017; // @[Mux.scala 31:69:@41222.4]
  wire [15:0] _T_97018; // @[Mux.scala 31:69:@41223.4]
  wire [15:0] _T_97019; // @[Mux.scala 31:69:@41224.4]
  wire [15:0] _T_97020; // @[Mux.scala 31:69:@41225.4]
  wire [15:0] _T_97021; // @[Mux.scala 31:69:@41226.4]
  wire [15:0] _T_97022; // @[Mux.scala 31:69:@41227.4]
  wire [15:0] _T_97023; // @[Mux.scala 31:69:@41228.4]
  wire [15:0] _T_97024; // @[Mux.scala 31:69:@41229.4]
  wire [15:0] _T_97025; // @[Mux.scala 31:69:@41230.4]
  wire [15:0] _T_97026; // @[Mux.scala 31:69:@41231.4]
  wire [15:0] _T_97027; // @[Mux.scala 31:69:@41232.4]
  wire [15:0] _T_97028; // @[Mux.scala 31:69:@41233.4]
  wire [15:0] _T_97029; // @[Mux.scala 31:69:@41234.4]
  wire  _T_97030; // @[OneHot.scala 66:30:@41235.4]
  wire  _T_97031; // @[OneHot.scala 66:30:@41236.4]
  wire  _T_97032; // @[OneHot.scala 66:30:@41237.4]
  wire  _T_97033; // @[OneHot.scala 66:30:@41238.4]
  wire  _T_97034; // @[OneHot.scala 66:30:@41239.4]
  wire  _T_97035; // @[OneHot.scala 66:30:@41240.4]
  wire  _T_97036; // @[OneHot.scala 66:30:@41241.4]
  wire  _T_97037; // @[OneHot.scala 66:30:@41242.4]
  wire  _T_97038; // @[OneHot.scala 66:30:@41243.4]
  wire  _T_97039; // @[OneHot.scala 66:30:@41244.4]
  wire  _T_97040; // @[OneHot.scala 66:30:@41245.4]
  wire  _T_97041; // @[OneHot.scala 66:30:@41246.4]
  wire  _T_97042; // @[OneHot.scala 66:30:@41247.4]
  wire  _T_97043; // @[OneHot.scala 66:30:@41248.4]
  wire  _T_97044; // @[OneHot.scala 66:30:@41249.4]
  wire  _T_97045; // @[OneHot.scala 66:30:@41250.4]
  wire [15:0] _T_97086; // @[Mux.scala 31:69:@41268.4]
  wire [15:0] _T_97087; // @[Mux.scala 31:69:@41269.4]
  wire [15:0] _T_97088; // @[Mux.scala 31:69:@41270.4]
  wire [15:0] _T_97089; // @[Mux.scala 31:69:@41271.4]
  wire [15:0] _T_97090; // @[Mux.scala 31:69:@41272.4]
  wire [15:0] _T_97091; // @[Mux.scala 31:69:@41273.4]
  wire [15:0] _T_97092; // @[Mux.scala 31:69:@41274.4]
  wire [15:0] _T_97093; // @[Mux.scala 31:69:@41275.4]
  wire [15:0] _T_97094; // @[Mux.scala 31:69:@41276.4]
  wire [15:0] _T_97095; // @[Mux.scala 31:69:@41277.4]
  wire [15:0] _T_97096; // @[Mux.scala 31:69:@41278.4]
  wire [15:0] _T_97097; // @[Mux.scala 31:69:@41279.4]
  wire [15:0] _T_97098; // @[Mux.scala 31:69:@41280.4]
  wire [15:0] _T_97099; // @[Mux.scala 31:69:@41281.4]
  wire [15:0] _T_97100; // @[Mux.scala 31:69:@41282.4]
  wire [15:0] _T_97101; // @[Mux.scala 31:69:@41283.4]
  wire  _T_97102; // @[OneHot.scala 66:30:@41284.4]
  wire  _T_97103; // @[OneHot.scala 66:30:@41285.4]
  wire  _T_97104; // @[OneHot.scala 66:30:@41286.4]
  wire  _T_97105; // @[OneHot.scala 66:30:@41287.4]
  wire  _T_97106; // @[OneHot.scala 66:30:@41288.4]
  wire  _T_97107; // @[OneHot.scala 66:30:@41289.4]
  wire  _T_97108; // @[OneHot.scala 66:30:@41290.4]
  wire  _T_97109; // @[OneHot.scala 66:30:@41291.4]
  wire  _T_97110; // @[OneHot.scala 66:30:@41292.4]
  wire  _T_97111; // @[OneHot.scala 66:30:@41293.4]
  wire  _T_97112; // @[OneHot.scala 66:30:@41294.4]
  wire  _T_97113; // @[OneHot.scala 66:30:@41295.4]
  wire  _T_97114; // @[OneHot.scala 66:30:@41296.4]
  wire  _T_97115; // @[OneHot.scala 66:30:@41297.4]
  wire  _T_97116; // @[OneHot.scala 66:30:@41298.4]
  wire  _T_97117; // @[OneHot.scala 66:30:@41299.4]
  wire [15:0] _T_97158; // @[Mux.scala 31:69:@41317.4]
  wire [15:0] _T_97159; // @[Mux.scala 31:69:@41318.4]
  wire [15:0] _T_97160; // @[Mux.scala 31:69:@41319.4]
  wire [15:0] _T_97161; // @[Mux.scala 31:69:@41320.4]
  wire [15:0] _T_97162; // @[Mux.scala 31:69:@41321.4]
  wire [15:0] _T_97163; // @[Mux.scala 31:69:@41322.4]
  wire [15:0] _T_97164; // @[Mux.scala 31:69:@41323.4]
  wire [15:0] _T_97165; // @[Mux.scala 31:69:@41324.4]
  wire [15:0] _T_97166; // @[Mux.scala 31:69:@41325.4]
  wire [15:0] _T_97167; // @[Mux.scala 31:69:@41326.4]
  wire [15:0] _T_97168; // @[Mux.scala 31:69:@41327.4]
  wire [15:0] _T_97169; // @[Mux.scala 31:69:@41328.4]
  wire [15:0] _T_97170; // @[Mux.scala 31:69:@41329.4]
  wire [15:0] _T_97171; // @[Mux.scala 31:69:@41330.4]
  wire [15:0] _T_97172; // @[Mux.scala 31:69:@41331.4]
  wire [15:0] _T_97173; // @[Mux.scala 31:69:@41332.4]
  wire  _T_97174; // @[OneHot.scala 66:30:@41333.4]
  wire  _T_97175; // @[OneHot.scala 66:30:@41334.4]
  wire  _T_97176; // @[OneHot.scala 66:30:@41335.4]
  wire  _T_97177; // @[OneHot.scala 66:30:@41336.4]
  wire  _T_97178; // @[OneHot.scala 66:30:@41337.4]
  wire  _T_97179; // @[OneHot.scala 66:30:@41338.4]
  wire  _T_97180; // @[OneHot.scala 66:30:@41339.4]
  wire  _T_97181; // @[OneHot.scala 66:30:@41340.4]
  wire  _T_97182; // @[OneHot.scala 66:30:@41341.4]
  wire  _T_97183; // @[OneHot.scala 66:30:@41342.4]
  wire  _T_97184; // @[OneHot.scala 66:30:@41343.4]
  wire  _T_97185; // @[OneHot.scala 66:30:@41344.4]
  wire  _T_97186; // @[OneHot.scala 66:30:@41345.4]
  wire  _T_97187; // @[OneHot.scala 66:30:@41346.4]
  wire  _T_97188; // @[OneHot.scala 66:30:@41347.4]
  wire  _T_97189; // @[OneHot.scala 66:30:@41348.4]
  wire [15:0] _T_97230; // @[Mux.scala 31:69:@41366.4]
  wire [15:0] _T_97231; // @[Mux.scala 31:69:@41367.4]
  wire [15:0] _T_97232; // @[Mux.scala 31:69:@41368.4]
  wire [15:0] _T_97233; // @[Mux.scala 31:69:@41369.4]
  wire [15:0] _T_97234; // @[Mux.scala 31:69:@41370.4]
  wire [15:0] _T_97235; // @[Mux.scala 31:69:@41371.4]
  wire [15:0] _T_97236; // @[Mux.scala 31:69:@41372.4]
  wire [15:0] _T_97237; // @[Mux.scala 31:69:@41373.4]
  wire [15:0] _T_97238; // @[Mux.scala 31:69:@41374.4]
  wire [15:0] _T_97239; // @[Mux.scala 31:69:@41375.4]
  wire [15:0] _T_97240; // @[Mux.scala 31:69:@41376.4]
  wire [15:0] _T_97241; // @[Mux.scala 31:69:@41377.4]
  wire [15:0] _T_97242; // @[Mux.scala 31:69:@41378.4]
  wire [15:0] _T_97243; // @[Mux.scala 31:69:@41379.4]
  wire [15:0] _T_97244; // @[Mux.scala 31:69:@41380.4]
  wire [15:0] _T_97245; // @[Mux.scala 31:69:@41381.4]
  wire  _T_97246; // @[OneHot.scala 66:30:@41382.4]
  wire  _T_97247; // @[OneHot.scala 66:30:@41383.4]
  wire  _T_97248; // @[OneHot.scala 66:30:@41384.4]
  wire  _T_97249; // @[OneHot.scala 66:30:@41385.4]
  wire  _T_97250; // @[OneHot.scala 66:30:@41386.4]
  wire  _T_97251; // @[OneHot.scala 66:30:@41387.4]
  wire  _T_97252; // @[OneHot.scala 66:30:@41388.4]
  wire  _T_97253; // @[OneHot.scala 66:30:@41389.4]
  wire  _T_97254; // @[OneHot.scala 66:30:@41390.4]
  wire  _T_97255; // @[OneHot.scala 66:30:@41391.4]
  wire  _T_97256; // @[OneHot.scala 66:30:@41392.4]
  wire  _T_97257; // @[OneHot.scala 66:30:@41393.4]
  wire  _T_97258; // @[OneHot.scala 66:30:@41394.4]
  wire  _T_97259; // @[OneHot.scala 66:30:@41395.4]
  wire  _T_97260; // @[OneHot.scala 66:30:@41396.4]
  wire  _T_97261; // @[OneHot.scala 66:30:@41397.4]
  wire [15:0] _T_97302; // @[Mux.scala 31:69:@41415.4]
  wire [15:0] _T_97303; // @[Mux.scala 31:69:@41416.4]
  wire [15:0] _T_97304; // @[Mux.scala 31:69:@41417.4]
  wire [15:0] _T_97305; // @[Mux.scala 31:69:@41418.4]
  wire [15:0] _T_97306; // @[Mux.scala 31:69:@41419.4]
  wire [15:0] _T_97307; // @[Mux.scala 31:69:@41420.4]
  wire [15:0] _T_97308; // @[Mux.scala 31:69:@41421.4]
  wire [15:0] _T_97309; // @[Mux.scala 31:69:@41422.4]
  wire [15:0] _T_97310; // @[Mux.scala 31:69:@41423.4]
  wire [15:0] _T_97311; // @[Mux.scala 31:69:@41424.4]
  wire [15:0] _T_97312; // @[Mux.scala 31:69:@41425.4]
  wire [15:0] _T_97313; // @[Mux.scala 31:69:@41426.4]
  wire [15:0] _T_97314; // @[Mux.scala 31:69:@41427.4]
  wire [15:0] _T_97315; // @[Mux.scala 31:69:@41428.4]
  wire [15:0] _T_97316; // @[Mux.scala 31:69:@41429.4]
  wire [15:0] _T_97317; // @[Mux.scala 31:69:@41430.4]
  wire  _T_97318; // @[OneHot.scala 66:30:@41431.4]
  wire  _T_97319; // @[OneHot.scala 66:30:@41432.4]
  wire  _T_97320; // @[OneHot.scala 66:30:@41433.4]
  wire  _T_97321; // @[OneHot.scala 66:30:@41434.4]
  wire  _T_97322; // @[OneHot.scala 66:30:@41435.4]
  wire  _T_97323; // @[OneHot.scala 66:30:@41436.4]
  wire  _T_97324; // @[OneHot.scala 66:30:@41437.4]
  wire  _T_97325; // @[OneHot.scala 66:30:@41438.4]
  wire  _T_97326; // @[OneHot.scala 66:30:@41439.4]
  wire  _T_97327; // @[OneHot.scala 66:30:@41440.4]
  wire  _T_97328; // @[OneHot.scala 66:30:@41441.4]
  wire  _T_97329; // @[OneHot.scala 66:30:@41442.4]
  wire  _T_97330; // @[OneHot.scala 66:30:@41443.4]
  wire  _T_97331; // @[OneHot.scala 66:30:@41444.4]
  wire  _T_97332; // @[OneHot.scala 66:30:@41445.4]
  wire  _T_97333; // @[OneHot.scala 66:30:@41446.4]
  wire [7:0] _T_97398; // @[Mux.scala 19:72:@41470.4]
  wire [15:0] _T_97406; // @[Mux.scala 19:72:@41478.4]
  wire [15:0] _T_97408; // @[Mux.scala 19:72:@41479.4]
  wire [7:0] _T_97415; // @[Mux.scala 19:72:@41486.4]
  wire [15:0] _T_97423; // @[Mux.scala 19:72:@41494.4]
  wire [15:0] _T_97425; // @[Mux.scala 19:72:@41495.4]
  wire [7:0] _T_97432; // @[Mux.scala 19:72:@41502.4]
  wire [15:0] _T_97440; // @[Mux.scala 19:72:@41510.4]
  wire [15:0] _T_97442; // @[Mux.scala 19:72:@41511.4]
  wire [7:0] _T_97449; // @[Mux.scala 19:72:@41518.4]
  wire [15:0] _T_97457; // @[Mux.scala 19:72:@41526.4]
  wire [15:0] _T_97459; // @[Mux.scala 19:72:@41527.4]
  wire [7:0] _T_97466; // @[Mux.scala 19:72:@41534.4]
  wire [15:0] _T_97474; // @[Mux.scala 19:72:@41542.4]
  wire [15:0] _T_97476; // @[Mux.scala 19:72:@41543.4]
  wire [7:0] _T_97483; // @[Mux.scala 19:72:@41550.4]
  wire [15:0] _T_97491; // @[Mux.scala 19:72:@41558.4]
  wire [15:0] _T_97493; // @[Mux.scala 19:72:@41559.4]
  wire [7:0] _T_97500; // @[Mux.scala 19:72:@41566.4]
  wire [15:0] _T_97508; // @[Mux.scala 19:72:@41574.4]
  wire [15:0] _T_97510; // @[Mux.scala 19:72:@41575.4]
  wire [7:0] _T_97517; // @[Mux.scala 19:72:@41582.4]
  wire [15:0] _T_97525; // @[Mux.scala 19:72:@41590.4]
  wire [15:0] _T_97527; // @[Mux.scala 19:72:@41591.4]
  wire [7:0] _T_97534; // @[Mux.scala 19:72:@41598.4]
  wire [15:0] _T_97542; // @[Mux.scala 19:72:@41606.4]
  wire [15:0] _T_97544; // @[Mux.scala 19:72:@41607.4]
  wire [7:0] _T_97551; // @[Mux.scala 19:72:@41614.4]
  wire [15:0] _T_97559; // @[Mux.scala 19:72:@41622.4]
  wire [15:0] _T_97561; // @[Mux.scala 19:72:@41623.4]
  wire [7:0] _T_97568; // @[Mux.scala 19:72:@41630.4]
  wire [15:0] _T_97576; // @[Mux.scala 19:72:@41638.4]
  wire [15:0] _T_97578; // @[Mux.scala 19:72:@41639.4]
  wire [7:0] _T_97585; // @[Mux.scala 19:72:@41646.4]
  wire [15:0] _T_97593; // @[Mux.scala 19:72:@41654.4]
  wire [15:0] _T_97595; // @[Mux.scala 19:72:@41655.4]
  wire [7:0] _T_97602; // @[Mux.scala 19:72:@41662.4]
  wire [15:0] _T_97610; // @[Mux.scala 19:72:@41670.4]
  wire [15:0] _T_97612; // @[Mux.scala 19:72:@41671.4]
  wire [7:0] _T_97619; // @[Mux.scala 19:72:@41678.4]
  wire [15:0] _T_97627; // @[Mux.scala 19:72:@41686.4]
  wire [15:0] _T_97629; // @[Mux.scala 19:72:@41687.4]
  wire [7:0] _T_97636; // @[Mux.scala 19:72:@41694.4]
  wire [15:0] _T_97644; // @[Mux.scala 19:72:@41702.4]
  wire [15:0] _T_97646; // @[Mux.scala 19:72:@41703.4]
  wire [7:0] _T_97653; // @[Mux.scala 19:72:@41710.4]
  wire [15:0] _T_97661; // @[Mux.scala 19:72:@41718.4]
  wire [15:0] _T_97663; // @[Mux.scala 19:72:@41719.4]
  wire [15:0] _T_97664; // @[Mux.scala 19:72:@41720.4]
  wire [15:0] _T_97665; // @[Mux.scala 19:72:@41721.4]
  wire [15:0] _T_97666; // @[Mux.scala 19:72:@41722.4]
  wire [15:0] _T_97667; // @[Mux.scala 19:72:@41723.4]
  wire [15:0] _T_97668; // @[Mux.scala 19:72:@41724.4]
  wire [15:0] _T_97669; // @[Mux.scala 19:72:@41725.4]
  wire [15:0] _T_97670; // @[Mux.scala 19:72:@41726.4]
  wire [15:0] _T_97671; // @[Mux.scala 19:72:@41727.4]
  wire [15:0] _T_97672; // @[Mux.scala 19:72:@41728.4]
  wire [15:0] _T_97673; // @[Mux.scala 19:72:@41729.4]
  wire [15:0] _T_97674; // @[Mux.scala 19:72:@41730.4]
  wire [15:0] _T_97675; // @[Mux.scala 19:72:@41731.4]
  wire [15:0] _T_97676; // @[Mux.scala 19:72:@41732.4]
  wire [15:0] _T_97677; // @[Mux.scala 19:72:@41733.4]
  wire [15:0] _T_97678; // @[Mux.scala 19:72:@41734.4]
  wire  outputPriorityPorts_0_0; // @[Mux.scala 19:72:@41738.4]
  wire  outputPriorityPorts_0_1; // @[Mux.scala 19:72:@41740.4]
  wire  outputPriorityPorts_0_2; // @[Mux.scala 19:72:@41742.4]
  wire  outputPriorityPorts_0_3; // @[Mux.scala 19:72:@41744.4]
  wire  outputPriorityPorts_0_4; // @[Mux.scala 19:72:@41746.4]
  wire  outputPriorityPorts_0_5; // @[Mux.scala 19:72:@41748.4]
  wire  outputPriorityPorts_0_6; // @[Mux.scala 19:72:@41750.4]
  wire  outputPriorityPorts_0_7; // @[Mux.scala 19:72:@41752.4]
  wire  outputPriorityPorts_0_8; // @[Mux.scala 19:72:@41754.4]
  wire  outputPriorityPorts_0_9; // @[Mux.scala 19:72:@41756.4]
  wire  outputPriorityPorts_0_10; // @[Mux.scala 19:72:@41758.4]
  wire  outputPriorityPorts_0_11; // @[Mux.scala 19:72:@41760.4]
  wire  outputPriorityPorts_0_12; // @[Mux.scala 19:72:@41762.4]
  wire  outputPriorityPorts_0_13; // @[Mux.scala 19:72:@41764.4]
  wire  outputPriorityPorts_0_14; // @[Mux.scala 19:72:@41766.4]
  wire  outputPriorityPorts_0_15; // @[Mux.scala 19:72:@41768.4]
  wire  _T_97822; // @[LoadQueue.scala 298:83:@41787.4]
  wire  _T_97825; // @[LoadQueue.scala 298:83:@41789.4]
  wire  _T_97828; // @[LoadQueue.scala 298:83:@41791.4]
  wire  _T_97831; // @[LoadQueue.scala 298:83:@41793.4]
  wire  _T_97834; // @[LoadQueue.scala 298:83:@41795.4]
  wire  _T_97837; // @[LoadQueue.scala 298:83:@41797.4]
  wire  _T_97840; // @[LoadQueue.scala 298:83:@41799.4]
  wire  _T_97843; // @[LoadQueue.scala 298:83:@41801.4]
  wire  _T_97846; // @[LoadQueue.scala 298:83:@41803.4]
  wire  _T_97849; // @[LoadQueue.scala 298:83:@41805.4]
  wire  _T_97852; // @[LoadQueue.scala 298:83:@41807.4]
  wire  _T_97855; // @[LoadQueue.scala 298:83:@41809.4]
  wire  _T_97858; // @[LoadQueue.scala 298:83:@41811.4]
  wire  _T_97861; // @[LoadQueue.scala 298:83:@41813.4]
  wire  _T_97864; // @[LoadQueue.scala 298:83:@41815.4]
  wire  _T_97867; // @[LoadQueue.scala 298:83:@41817.4]
  wire [15:0] _T_97950; // @[Mux.scala 31:69:@41871.4]
  wire [15:0] _T_97951; // @[Mux.scala 31:69:@41872.4]
  wire [15:0] _T_97952; // @[Mux.scala 31:69:@41873.4]
  wire [15:0] _T_97953; // @[Mux.scala 31:69:@41874.4]
  wire [15:0] _T_97954; // @[Mux.scala 31:69:@41875.4]
  wire [15:0] _T_97955; // @[Mux.scala 31:69:@41876.4]
  wire [15:0] _T_97956; // @[Mux.scala 31:69:@41877.4]
  wire [15:0] _T_97957; // @[Mux.scala 31:69:@41878.4]
  wire [15:0] _T_97958; // @[Mux.scala 31:69:@41879.4]
  wire [15:0] _T_97959; // @[Mux.scala 31:69:@41880.4]
  wire [15:0] _T_97960; // @[Mux.scala 31:69:@41881.4]
  wire [15:0] _T_97961; // @[Mux.scala 31:69:@41882.4]
  wire [15:0] _T_97962; // @[Mux.scala 31:69:@41883.4]
  wire [15:0] _T_97963; // @[Mux.scala 31:69:@41884.4]
  wire [15:0] _T_97964; // @[Mux.scala 31:69:@41885.4]
  wire [15:0] _T_97965; // @[Mux.scala 31:69:@41886.4]
  wire  _T_97966; // @[OneHot.scala 66:30:@41887.4]
  wire  _T_97967; // @[OneHot.scala 66:30:@41888.4]
  wire  _T_97968; // @[OneHot.scala 66:30:@41889.4]
  wire  _T_97969; // @[OneHot.scala 66:30:@41890.4]
  wire  _T_97970; // @[OneHot.scala 66:30:@41891.4]
  wire  _T_97971; // @[OneHot.scala 66:30:@41892.4]
  wire  _T_97972; // @[OneHot.scala 66:30:@41893.4]
  wire  _T_97973; // @[OneHot.scala 66:30:@41894.4]
  wire  _T_97974; // @[OneHot.scala 66:30:@41895.4]
  wire  _T_97975; // @[OneHot.scala 66:30:@41896.4]
  wire  _T_97976; // @[OneHot.scala 66:30:@41897.4]
  wire  _T_97977; // @[OneHot.scala 66:30:@41898.4]
  wire  _T_97978; // @[OneHot.scala 66:30:@41899.4]
  wire  _T_97979; // @[OneHot.scala 66:30:@41900.4]
  wire  _T_97980; // @[OneHot.scala 66:30:@41901.4]
  wire  _T_97981; // @[OneHot.scala 66:30:@41902.4]
  wire [15:0] _T_98022; // @[Mux.scala 31:69:@41920.4]
  wire [15:0] _T_98023; // @[Mux.scala 31:69:@41921.4]
  wire [15:0] _T_98024; // @[Mux.scala 31:69:@41922.4]
  wire [15:0] _T_98025; // @[Mux.scala 31:69:@41923.4]
  wire [15:0] _T_98026; // @[Mux.scala 31:69:@41924.4]
  wire [15:0] _T_98027; // @[Mux.scala 31:69:@41925.4]
  wire [15:0] _T_98028; // @[Mux.scala 31:69:@41926.4]
  wire [15:0] _T_98029; // @[Mux.scala 31:69:@41927.4]
  wire [15:0] _T_98030; // @[Mux.scala 31:69:@41928.4]
  wire [15:0] _T_98031; // @[Mux.scala 31:69:@41929.4]
  wire [15:0] _T_98032; // @[Mux.scala 31:69:@41930.4]
  wire [15:0] _T_98033; // @[Mux.scala 31:69:@41931.4]
  wire [15:0] _T_98034; // @[Mux.scala 31:69:@41932.4]
  wire [15:0] _T_98035; // @[Mux.scala 31:69:@41933.4]
  wire [15:0] _T_98036; // @[Mux.scala 31:69:@41934.4]
  wire [15:0] _T_98037; // @[Mux.scala 31:69:@41935.4]
  wire  _T_98038; // @[OneHot.scala 66:30:@41936.4]
  wire  _T_98039; // @[OneHot.scala 66:30:@41937.4]
  wire  _T_98040; // @[OneHot.scala 66:30:@41938.4]
  wire  _T_98041; // @[OneHot.scala 66:30:@41939.4]
  wire  _T_98042; // @[OneHot.scala 66:30:@41940.4]
  wire  _T_98043; // @[OneHot.scala 66:30:@41941.4]
  wire  _T_98044; // @[OneHot.scala 66:30:@41942.4]
  wire  _T_98045; // @[OneHot.scala 66:30:@41943.4]
  wire  _T_98046; // @[OneHot.scala 66:30:@41944.4]
  wire  _T_98047; // @[OneHot.scala 66:30:@41945.4]
  wire  _T_98048; // @[OneHot.scala 66:30:@41946.4]
  wire  _T_98049; // @[OneHot.scala 66:30:@41947.4]
  wire  _T_98050; // @[OneHot.scala 66:30:@41948.4]
  wire  _T_98051; // @[OneHot.scala 66:30:@41949.4]
  wire  _T_98052; // @[OneHot.scala 66:30:@41950.4]
  wire  _T_98053; // @[OneHot.scala 66:30:@41951.4]
  wire [15:0] _T_98094; // @[Mux.scala 31:69:@41969.4]
  wire [15:0] _T_98095; // @[Mux.scala 31:69:@41970.4]
  wire [15:0] _T_98096; // @[Mux.scala 31:69:@41971.4]
  wire [15:0] _T_98097; // @[Mux.scala 31:69:@41972.4]
  wire [15:0] _T_98098; // @[Mux.scala 31:69:@41973.4]
  wire [15:0] _T_98099; // @[Mux.scala 31:69:@41974.4]
  wire [15:0] _T_98100; // @[Mux.scala 31:69:@41975.4]
  wire [15:0] _T_98101; // @[Mux.scala 31:69:@41976.4]
  wire [15:0] _T_98102; // @[Mux.scala 31:69:@41977.4]
  wire [15:0] _T_98103; // @[Mux.scala 31:69:@41978.4]
  wire [15:0] _T_98104; // @[Mux.scala 31:69:@41979.4]
  wire [15:0] _T_98105; // @[Mux.scala 31:69:@41980.4]
  wire [15:0] _T_98106; // @[Mux.scala 31:69:@41981.4]
  wire [15:0] _T_98107; // @[Mux.scala 31:69:@41982.4]
  wire [15:0] _T_98108; // @[Mux.scala 31:69:@41983.4]
  wire [15:0] _T_98109; // @[Mux.scala 31:69:@41984.4]
  wire  _T_98110; // @[OneHot.scala 66:30:@41985.4]
  wire  _T_98111; // @[OneHot.scala 66:30:@41986.4]
  wire  _T_98112; // @[OneHot.scala 66:30:@41987.4]
  wire  _T_98113; // @[OneHot.scala 66:30:@41988.4]
  wire  _T_98114; // @[OneHot.scala 66:30:@41989.4]
  wire  _T_98115; // @[OneHot.scala 66:30:@41990.4]
  wire  _T_98116; // @[OneHot.scala 66:30:@41991.4]
  wire  _T_98117; // @[OneHot.scala 66:30:@41992.4]
  wire  _T_98118; // @[OneHot.scala 66:30:@41993.4]
  wire  _T_98119; // @[OneHot.scala 66:30:@41994.4]
  wire  _T_98120; // @[OneHot.scala 66:30:@41995.4]
  wire  _T_98121; // @[OneHot.scala 66:30:@41996.4]
  wire  _T_98122; // @[OneHot.scala 66:30:@41997.4]
  wire  _T_98123; // @[OneHot.scala 66:30:@41998.4]
  wire  _T_98124; // @[OneHot.scala 66:30:@41999.4]
  wire  _T_98125; // @[OneHot.scala 66:30:@42000.4]
  wire [15:0] _T_98166; // @[Mux.scala 31:69:@42018.4]
  wire [15:0] _T_98167; // @[Mux.scala 31:69:@42019.4]
  wire [15:0] _T_98168; // @[Mux.scala 31:69:@42020.4]
  wire [15:0] _T_98169; // @[Mux.scala 31:69:@42021.4]
  wire [15:0] _T_98170; // @[Mux.scala 31:69:@42022.4]
  wire [15:0] _T_98171; // @[Mux.scala 31:69:@42023.4]
  wire [15:0] _T_98172; // @[Mux.scala 31:69:@42024.4]
  wire [15:0] _T_98173; // @[Mux.scala 31:69:@42025.4]
  wire [15:0] _T_98174; // @[Mux.scala 31:69:@42026.4]
  wire [15:0] _T_98175; // @[Mux.scala 31:69:@42027.4]
  wire [15:0] _T_98176; // @[Mux.scala 31:69:@42028.4]
  wire [15:0] _T_98177; // @[Mux.scala 31:69:@42029.4]
  wire [15:0] _T_98178; // @[Mux.scala 31:69:@42030.4]
  wire [15:0] _T_98179; // @[Mux.scala 31:69:@42031.4]
  wire [15:0] _T_98180; // @[Mux.scala 31:69:@42032.4]
  wire [15:0] _T_98181; // @[Mux.scala 31:69:@42033.4]
  wire  _T_98182; // @[OneHot.scala 66:30:@42034.4]
  wire  _T_98183; // @[OneHot.scala 66:30:@42035.4]
  wire  _T_98184; // @[OneHot.scala 66:30:@42036.4]
  wire  _T_98185; // @[OneHot.scala 66:30:@42037.4]
  wire  _T_98186; // @[OneHot.scala 66:30:@42038.4]
  wire  _T_98187; // @[OneHot.scala 66:30:@42039.4]
  wire  _T_98188; // @[OneHot.scala 66:30:@42040.4]
  wire  _T_98189; // @[OneHot.scala 66:30:@42041.4]
  wire  _T_98190; // @[OneHot.scala 66:30:@42042.4]
  wire  _T_98191; // @[OneHot.scala 66:30:@42043.4]
  wire  _T_98192; // @[OneHot.scala 66:30:@42044.4]
  wire  _T_98193; // @[OneHot.scala 66:30:@42045.4]
  wire  _T_98194; // @[OneHot.scala 66:30:@42046.4]
  wire  _T_98195; // @[OneHot.scala 66:30:@42047.4]
  wire  _T_98196; // @[OneHot.scala 66:30:@42048.4]
  wire  _T_98197; // @[OneHot.scala 66:30:@42049.4]
  wire [15:0] _T_98238; // @[Mux.scala 31:69:@42067.4]
  wire [15:0] _T_98239; // @[Mux.scala 31:69:@42068.4]
  wire [15:0] _T_98240; // @[Mux.scala 31:69:@42069.4]
  wire [15:0] _T_98241; // @[Mux.scala 31:69:@42070.4]
  wire [15:0] _T_98242; // @[Mux.scala 31:69:@42071.4]
  wire [15:0] _T_98243; // @[Mux.scala 31:69:@42072.4]
  wire [15:0] _T_98244; // @[Mux.scala 31:69:@42073.4]
  wire [15:0] _T_98245; // @[Mux.scala 31:69:@42074.4]
  wire [15:0] _T_98246; // @[Mux.scala 31:69:@42075.4]
  wire [15:0] _T_98247; // @[Mux.scala 31:69:@42076.4]
  wire [15:0] _T_98248; // @[Mux.scala 31:69:@42077.4]
  wire [15:0] _T_98249; // @[Mux.scala 31:69:@42078.4]
  wire [15:0] _T_98250; // @[Mux.scala 31:69:@42079.4]
  wire [15:0] _T_98251; // @[Mux.scala 31:69:@42080.4]
  wire [15:0] _T_98252; // @[Mux.scala 31:69:@42081.4]
  wire [15:0] _T_98253; // @[Mux.scala 31:69:@42082.4]
  wire  _T_98254; // @[OneHot.scala 66:30:@42083.4]
  wire  _T_98255; // @[OneHot.scala 66:30:@42084.4]
  wire  _T_98256; // @[OneHot.scala 66:30:@42085.4]
  wire  _T_98257; // @[OneHot.scala 66:30:@42086.4]
  wire  _T_98258; // @[OneHot.scala 66:30:@42087.4]
  wire  _T_98259; // @[OneHot.scala 66:30:@42088.4]
  wire  _T_98260; // @[OneHot.scala 66:30:@42089.4]
  wire  _T_98261; // @[OneHot.scala 66:30:@42090.4]
  wire  _T_98262; // @[OneHot.scala 66:30:@42091.4]
  wire  _T_98263; // @[OneHot.scala 66:30:@42092.4]
  wire  _T_98264; // @[OneHot.scala 66:30:@42093.4]
  wire  _T_98265; // @[OneHot.scala 66:30:@42094.4]
  wire  _T_98266; // @[OneHot.scala 66:30:@42095.4]
  wire  _T_98267; // @[OneHot.scala 66:30:@42096.4]
  wire  _T_98268; // @[OneHot.scala 66:30:@42097.4]
  wire  _T_98269; // @[OneHot.scala 66:30:@42098.4]
  wire [15:0] _T_98310; // @[Mux.scala 31:69:@42116.4]
  wire [15:0] _T_98311; // @[Mux.scala 31:69:@42117.4]
  wire [15:0] _T_98312; // @[Mux.scala 31:69:@42118.4]
  wire [15:0] _T_98313; // @[Mux.scala 31:69:@42119.4]
  wire [15:0] _T_98314; // @[Mux.scala 31:69:@42120.4]
  wire [15:0] _T_98315; // @[Mux.scala 31:69:@42121.4]
  wire [15:0] _T_98316; // @[Mux.scala 31:69:@42122.4]
  wire [15:0] _T_98317; // @[Mux.scala 31:69:@42123.4]
  wire [15:0] _T_98318; // @[Mux.scala 31:69:@42124.4]
  wire [15:0] _T_98319; // @[Mux.scala 31:69:@42125.4]
  wire [15:0] _T_98320; // @[Mux.scala 31:69:@42126.4]
  wire [15:0] _T_98321; // @[Mux.scala 31:69:@42127.4]
  wire [15:0] _T_98322; // @[Mux.scala 31:69:@42128.4]
  wire [15:0] _T_98323; // @[Mux.scala 31:69:@42129.4]
  wire [15:0] _T_98324; // @[Mux.scala 31:69:@42130.4]
  wire [15:0] _T_98325; // @[Mux.scala 31:69:@42131.4]
  wire  _T_98326; // @[OneHot.scala 66:30:@42132.4]
  wire  _T_98327; // @[OneHot.scala 66:30:@42133.4]
  wire  _T_98328; // @[OneHot.scala 66:30:@42134.4]
  wire  _T_98329; // @[OneHot.scala 66:30:@42135.4]
  wire  _T_98330; // @[OneHot.scala 66:30:@42136.4]
  wire  _T_98331; // @[OneHot.scala 66:30:@42137.4]
  wire  _T_98332; // @[OneHot.scala 66:30:@42138.4]
  wire  _T_98333; // @[OneHot.scala 66:30:@42139.4]
  wire  _T_98334; // @[OneHot.scala 66:30:@42140.4]
  wire  _T_98335; // @[OneHot.scala 66:30:@42141.4]
  wire  _T_98336; // @[OneHot.scala 66:30:@42142.4]
  wire  _T_98337; // @[OneHot.scala 66:30:@42143.4]
  wire  _T_98338; // @[OneHot.scala 66:30:@42144.4]
  wire  _T_98339; // @[OneHot.scala 66:30:@42145.4]
  wire  _T_98340; // @[OneHot.scala 66:30:@42146.4]
  wire  _T_98341; // @[OneHot.scala 66:30:@42147.4]
  wire [15:0] _T_98382; // @[Mux.scala 31:69:@42165.4]
  wire [15:0] _T_98383; // @[Mux.scala 31:69:@42166.4]
  wire [15:0] _T_98384; // @[Mux.scala 31:69:@42167.4]
  wire [15:0] _T_98385; // @[Mux.scala 31:69:@42168.4]
  wire [15:0] _T_98386; // @[Mux.scala 31:69:@42169.4]
  wire [15:0] _T_98387; // @[Mux.scala 31:69:@42170.4]
  wire [15:0] _T_98388; // @[Mux.scala 31:69:@42171.4]
  wire [15:0] _T_98389; // @[Mux.scala 31:69:@42172.4]
  wire [15:0] _T_98390; // @[Mux.scala 31:69:@42173.4]
  wire [15:0] _T_98391; // @[Mux.scala 31:69:@42174.4]
  wire [15:0] _T_98392; // @[Mux.scala 31:69:@42175.4]
  wire [15:0] _T_98393; // @[Mux.scala 31:69:@42176.4]
  wire [15:0] _T_98394; // @[Mux.scala 31:69:@42177.4]
  wire [15:0] _T_98395; // @[Mux.scala 31:69:@42178.4]
  wire [15:0] _T_98396; // @[Mux.scala 31:69:@42179.4]
  wire [15:0] _T_98397; // @[Mux.scala 31:69:@42180.4]
  wire  _T_98398; // @[OneHot.scala 66:30:@42181.4]
  wire  _T_98399; // @[OneHot.scala 66:30:@42182.4]
  wire  _T_98400; // @[OneHot.scala 66:30:@42183.4]
  wire  _T_98401; // @[OneHot.scala 66:30:@42184.4]
  wire  _T_98402; // @[OneHot.scala 66:30:@42185.4]
  wire  _T_98403; // @[OneHot.scala 66:30:@42186.4]
  wire  _T_98404; // @[OneHot.scala 66:30:@42187.4]
  wire  _T_98405; // @[OneHot.scala 66:30:@42188.4]
  wire  _T_98406; // @[OneHot.scala 66:30:@42189.4]
  wire  _T_98407; // @[OneHot.scala 66:30:@42190.4]
  wire  _T_98408; // @[OneHot.scala 66:30:@42191.4]
  wire  _T_98409; // @[OneHot.scala 66:30:@42192.4]
  wire  _T_98410; // @[OneHot.scala 66:30:@42193.4]
  wire  _T_98411; // @[OneHot.scala 66:30:@42194.4]
  wire  _T_98412; // @[OneHot.scala 66:30:@42195.4]
  wire  _T_98413; // @[OneHot.scala 66:30:@42196.4]
  wire [15:0] _T_98454; // @[Mux.scala 31:69:@42214.4]
  wire [15:0] _T_98455; // @[Mux.scala 31:69:@42215.4]
  wire [15:0] _T_98456; // @[Mux.scala 31:69:@42216.4]
  wire [15:0] _T_98457; // @[Mux.scala 31:69:@42217.4]
  wire [15:0] _T_98458; // @[Mux.scala 31:69:@42218.4]
  wire [15:0] _T_98459; // @[Mux.scala 31:69:@42219.4]
  wire [15:0] _T_98460; // @[Mux.scala 31:69:@42220.4]
  wire [15:0] _T_98461; // @[Mux.scala 31:69:@42221.4]
  wire [15:0] _T_98462; // @[Mux.scala 31:69:@42222.4]
  wire [15:0] _T_98463; // @[Mux.scala 31:69:@42223.4]
  wire [15:0] _T_98464; // @[Mux.scala 31:69:@42224.4]
  wire [15:0] _T_98465; // @[Mux.scala 31:69:@42225.4]
  wire [15:0] _T_98466; // @[Mux.scala 31:69:@42226.4]
  wire [15:0] _T_98467; // @[Mux.scala 31:69:@42227.4]
  wire [15:0] _T_98468; // @[Mux.scala 31:69:@42228.4]
  wire [15:0] _T_98469; // @[Mux.scala 31:69:@42229.4]
  wire  _T_98470; // @[OneHot.scala 66:30:@42230.4]
  wire  _T_98471; // @[OneHot.scala 66:30:@42231.4]
  wire  _T_98472; // @[OneHot.scala 66:30:@42232.4]
  wire  _T_98473; // @[OneHot.scala 66:30:@42233.4]
  wire  _T_98474; // @[OneHot.scala 66:30:@42234.4]
  wire  _T_98475; // @[OneHot.scala 66:30:@42235.4]
  wire  _T_98476; // @[OneHot.scala 66:30:@42236.4]
  wire  _T_98477; // @[OneHot.scala 66:30:@42237.4]
  wire  _T_98478; // @[OneHot.scala 66:30:@42238.4]
  wire  _T_98479; // @[OneHot.scala 66:30:@42239.4]
  wire  _T_98480; // @[OneHot.scala 66:30:@42240.4]
  wire  _T_98481; // @[OneHot.scala 66:30:@42241.4]
  wire  _T_98482; // @[OneHot.scala 66:30:@42242.4]
  wire  _T_98483; // @[OneHot.scala 66:30:@42243.4]
  wire  _T_98484; // @[OneHot.scala 66:30:@42244.4]
  wire  _T_98485; // @[OneHot.scala 66:30:@42245.4]
  wire [15:0] _T_98526; // @[Mux.scala 31:69:@42263.4]
  wire [15:0] _T_98527; // @[Mux.scala 31:69:@42264.4]
  wire [15:0] _T_98528; // @[Mux.scala 31:69:@42265.4]
  wire [15:0] _T_98529; // @[Mux.scala 31:69:@42266.4]
  wire [15:0] _T_98530; // @[Mux.scala 31:69:@42267.4]
  wire [15:0] _T_98531; // @[Mux.scala 31:69:@42268.4]
  wire [15:0] _T_98532; // @[Mux.scala 31:69:@42269.4]
  wire [15:0] _T_98533; // @[Mux.scala 31:69:@42270.4]
  wire [15:0] _T_98534; // @[Mux.scala 31:69:@42271.4]
  wire [15:0] _T_98535; // @[Mux.scala 31:69:@42272.4]
  wire [15:0] _T_98536; // @[Mux.scala 31:69:@42273.4]
  wire [15:0] _T_98537; // @[Mux.scala 31:69:@42274.4]
  wire [15:0] _T_98538; // @[Mux.scala 31:69:@42275.4]
  wire [15:0] _T_98539; // @[Mux.scala 31:69:@42276.4]
  wire [15:0] _T_98540; // @[Mux.scala 31:69:@42277.4]
  wire [15:0] _T_98541; // @[Mux.scala 31:69:@42278.4]
  wire  _T_98542; // @[OneHot.scala 66:30:@42279.4]
  wire  _T_98543; // @[OneHot.scala 66:30:@42280.4]
  wire  _T_98544; // @[OneHot.scala 66:30:@42281.4]
  wire  _T_98545; // @[OneHot.scala 66:30:@42282.4]
  wire  _T_98546; // @[OneHot.scala 66:30:@42283.4]
  wire  _T_98547; // @[OneHot.scala 66:30:@42284.4]
  wire  _T_98548; // @[OneHot.scala 66:30:@42285.4]
  wire  _T_98549; // @[OneHot.scala 66:30:@42286.4]
  wire  _T_98550; // @[OneHot.scala 66:30:@42287.4]
  wire  _T_98551; // @[OneHot.scala 66:30:@42288.4]
  wire  _T_98552; // @[OneHot.scala 66:30:@42289.4]
  wire  _T_98553; // @[OneHot.scala 66:30:@42290.4]
  wire  _T_98554; // @[OneHot.scala 66:30:@42291.4]
  wire  _T_98555; // @[OneHot.scala 66:30:@42292.4]
  wire  _T_98556; // @[OneHot.scala 66:30:@42293.4]
  wire  _T_98557; // @[OneHot.scala 66:30:@42294.4]
  wire [15:0] _T_98598; // @[Mux.scala 31:69:@42312.4]
  wire [15:0] _T_98599; // @[Mux.scala 31:69:@42313.4]
  wire [15:0] _T_98600; // @[Mux.scala 31:69:@42314.4]
  wire [15:0] _T_98601; // @[Mux.scala 31:69:@42315.4]
  wire [15:0] _T_98602; // @[Mux.scala 31:69:@42316.4]
  wire [15:0] _T_98603; // @[Mux.scala 31:69:@42317.4]
  wire [15:0] _T_98604; // @[Mux.scala 31:69:@42318.4]
  wire [15:0] _T_98605; // @[Mux.scala 31:69:@42319.4]
  wire [15:0] _T_98606; // @[Mux.scala 31:69:@42320.4]
  wire [15:0] _T_98607; // @[Mux.scala 31:69:@42321.4]
  wire [15:0] _T_98608; // @[Mux.scala 31:69:@42322.4]
  wire [15:0] _T_98609; // @[Mux.scala 31:69:@42323.4]
  wire [15:0] _T_98610; // @[Mux.scala 31:69:@42324.4]
  wire [15:0] _T_98611; // @[Mux.scala 31:69:@42325.4]
  wire [15:0] _T_98612; // @[Mux.scala 31:69:@42326.4]
  wire [15:0] _T_98613; // @[Mux.scala 31:69:@42327.4]
  wire  _T_98614; // @[OneHot.scala 66:30:@42328.4]
  wire  _T_98615; // @[OneHot.scala 66:30:@42329.4]
  wire  _T_98616; // @[OneHot.scala 66:30:@42330.4]
  wire  _T_98617; // @[OneHot.scala 66:30:@42331.4]
  wire  _T_98618; // @[OneHot.scala 66:30:@42332.4]
  wire  _T_98619; // @[OneHot.scala 66:30:@42333.4]
  wire  _T_98620; // @[OneHot.scala 66:30:@42334.4]
  wire  _T_98621; // @[OneHot.scala 66:30:@42335.4]
  wire  _T_98622; // @[OneHot.scala 66:30:@42336.4]
  wire  _T_98623; // @[OneHot.scala 66:30:@42337.4]
  wire  _T_98624; // @[OneHot.scala 66:30:@42338.4]
  wire  _T_98625; // @[OneHot.scala 66:30:@42339.4]
  wire  _T_98626; // @[OneHot.scala 66:30:@42340.4]
  wire  _T_98627; // @[OneHot.scala 66:30:@42341.4]
  wire  _T_98628; // @[OneHot.scala 66:30:@42342.4]
  wire  _T_98629; // @[OneHot.scala 66:30:@42343.4]
  wire [15:0] _T_98670; // @[Mux.scala 31:69:@42361.4]
  wire [15:0] _T_98671; // @[Mux.scala 31:69:@42362.4]
  wire [15:0] _T_98672; // @[Mux.scala 31:69:@42363.4]
  wire [15:0] _T_98673; // @[Mux.scala 31:69:@42364.4]
  wire [15:0] _T_98674; // @[Mux.scala 31:69:@42365.4]
  wire [15:0] _T_98675; // @[Mux.scala 31:69:@42366.4]
  wire [15:0] _T_98676; // @[Mux.scala 31:69:@42367.4]
  wire [15:0] _T_98677; // @[Mux.scala 31:69:@42368.4]
  wire [15:0] _T_98678; // @[Mux.scala 31:69:@42369.4]
  wire [15:0] _T_98679; // @[Mux.scala 31:69:@42370.4]
  wire [15:0] _T_98680; // @[Mux.scala 31:69:@42371.4]
  wire [15:0] _T_98681; // @[Mux.scala 31:69:@42372.4]
  wire [15:0] _T_98682; // @[Mux.scala 31:69:@42373.4]
  wire [15:0] _T_98683; // @[Mux.scala 31:69:@42374.4]
  wire [15:0] _T_98684; // @[Mux.scala 31:69:@42375.4]
  wire [15:0] _T_98685; // @[Mux.scala 31:69:@42376.4]
  wire  _T_98686; // @[OneHot.scala 66:30:@42377.4]
  wire  _T_98687; // @[OneHot.scala 66:30:@42378.4]
  wire  _T_98688; // @[OneHot.scala 66:30:@42379.4]
  wire  _T_98689; // @[OneHot.scala 66:30:@42380.4]
  wire  _T_98690; // @[OneHot.scala 66:30:@42381.4]
  wire  _T_98691; // @[OneHot.scala 66:30:@42382.4]
  wire  _T_98692; // @[OneHot.scala 66:30:@42383.4]
  wire  _T_98693; // @[OneHot.scala 66:30:@42384.4]
  wire  _T_98694; // @[OneHot.scala 66:30:@42385.4]
  wire  _T_98695; // @[OneHot.scala 66:30:@42386.4]
  wire  _T_98696; // @[OneHot.scala 66:30:@42387.4]
  wire  _T_98697; // @[OneHot.scala 66:30:@42388.4]
  wire  _T_98698; // @[OneHot.scala 66:30:@42389.4]
  wire  _T_98699; // @[OneHot.scala 66:30:@42390.4]
  wire  _T_98700; // @[OneHot.scala 66:30:@42391.4]
  wire  _T_98701; // @[OneHot.scala 66:30:@42392.4]
  wire [15:0] _T_98742; // @[Mux.scala 31:69:@42410.4]
  wire [15:0] _T_98743; // @[Mux.scala 31:69:@42411.4]
  wire [15:0] _T_98744; // @[Mux.scala 31:69:@42412.4]
  wire [15:0] _T_98745; // @[Mux.scala 31:69:@42413.4]
  wire [15:0] _T_98746; // @[Mux.scala 31:69:@42414.4]
  wire [15:0] _T_98747; // @[Mux.scala 31:69:@42415.4]
  wire [15:0] _T_98748; // @[Mux.scala 31:69:@42416.4]
  wire [15:0] _T_98749; // @[Mux.scala 31:69:@42417.4]
  wire [15:0] _T_98750; // @[Mux.scala 31:69:@42418.4]
  wire [15:0] _T_98751; // @[Mux.scala 31:69:@42419.4]
  wire [15:0] _T_98752; // @[Mux.scala 31:69:@42420.4]
  wire [15:0] _T_98753; // @[Mux.scala 31:69:@42421.4]
  wire [15:0] _T_98754; // @[Mux.scala 31:69:@42422.4]
  wire [15:0] _T_98755; // @[Mux.scala 31:69:@42423.4]
  wire [15:0] _T_98756; // @[Mux.scala 31:69:@42424.4]
  wire [15:0] _T_98757; // @[Mux.scala 31:69:@42425.4]
  wire  _T_98758; // @[OneHot.scala 66:30:@42426.4]
  wire  _T_98759; // @[OneHot.scala 66:30:@42427.4]
  wire  _T_98760; // @[OneHot.scala 66:30:@42428.4]
  wire  _T_98761; // @[OneHot.scala 66:30:@42429.4]
  wire  _T_98762; // @[OneHot.scala 66:30:@42430.4]
  wire  _T_98763; // @[OneHot.scala 66:30:@42431.4]
  wire  _T_98764; // @[OneHot.scala 66:30:@42432.4]
  wire  _T_98765; // @[OneHot.scala 66:30:@42433.4]
  wire  _T_98766; // @[OneHot.scala 66:30:@42434.4]
  wire  _T_98767; // @[OneHot.scala 66:30:@42435.4]
  wire  _T_98768; // @[OneHot.scala 66:30:@42436.4]
  wire  _T_98769; // @[OneHot.scala 66:30:@42437.4]
  wire  _T_98770; // @[OneHot.scala 66:30:@42438.4]
  wire  _T_98771; // @[OneHot.scala 66:30:@42439.4]
  wire  _T_98772; // @[OneHot.scala 66:30:@42440.4]
  wire  _T_98773; // @[OneHot.scala 66:30:@42441.4]
  wire [15:0] _T_98814; // @[Mux.scala 31:69:@42459.4]
  wire [15:0] _T_98815; // @[Mux.scala 31:69:@42460.4]
  wire [15:0] _T_98816; // @[Mux.scala 31:69:@42461.4]
  wire [15:0] _T_98817; // @[Mux.scala 31:69:@42462.4]
  wire [15:0] _T_98818; // @[Mux.scala 31:69:@42463.4]
  wire [15:0] _T_98819; // @[Mux.scala 31:69:@42464.4]
  wire [15:0] _T_98820; // @[Mux.scala 31:69:@42465.4]
  wire [15:0] _T_98821; // @[Mux.scala 31:69:@42466.4]
  wire [15:0] _T_98822; // @[Mux.scala 31:69:@42467.4]
  wire [15:0] _T_98823; // @[Mux.scala 31:69:@42468.4]
  wire [15:0] _T_98824; // @[Mux.scala 31:69:@42469.4]
  wire [15:0] _T_98825; // @[Mux.scala 31:69:@42470.4]
  wire [15:0] _T_98826; // @[Mux.scala 31:69:@42471.4]
  wire [15:0] _T_98827; // @[Mux.scala 31:69:@42472.4]
  wire [15:0] _T_98828; // @[Mux.scala 31:69:@42473.4]
  wire [15:0] _T_98829; // @[Mux.scala 31:69:@42474.4]
  wire  _T_98830; // @[OneHot.scala 66:30:@42475.4]
  wire  _T_98831; // @[OneHot.scala 66:30:@42476.4]
  wire  _T_98832; // @[OneHot.scala 66:30:@42477.4]
  wire  _T_98833; // @[OneHot.scala 66:30:@42478.4]
  wire  _T_98834; // @[OneHot.scala 66:30:@42479.4]
  wire  _T_98835; // @[OneHot.scala 66:30:@42480.4]
  wire  _T_98836; // @[OneHot.scala 66:30:@42481.4]
  wire  _T_98837; // @[OneHot.scala 66:30:@42482.4]
  wire  _T_98838; // @[OneHot.scala 66:30:@42483.4]
  wire  _T_98839; // @[OneHot.scala 66:30:@42484.4]
  wire  _T_98840; // @[OneHot.scala 66:30:@42485.4]
  wire  _T_98841; // @[OneHot.scala 66:30:@42486.4]
  wire  _T_98842; // @[OneHot.scala 66:30:@42487.4]
  wire  _T_98843; // @[OneHot.scala 66:30:@42488.4]
  wire  _T_98844; // @[OneHot.scala 66:30:@42489.4]
  wire  _T_98845; // @[OneHot.scala 66:30:@42490.4]
  wire [15:0] _T_98886; // @[Mux.scala 31:69:@42508.4]
  wire [15:0] _T_98887; // @[Mux.scala 31:69:@42509.4]
  wire [15:0] _T_98888; // @[Mux.scala 31:69:@42510.4]
  wire [15:0] _T_98889; // @[Mux.scala 31:69:@42511.4]
  wire [15:0] _T_98890; // @[Mux.scala 31:69:@42512.4]
  wire [15:0] _T_98891; // @[Mux.scala 31:69:@42513.4]
  wire [15:0] _T_98892; // @[Mux.scala 31:69:@42514.4]
  wire [15:0] _T_98893; // @[Mux.scala 31:69:@42515.4]
  wire [15:0] _T_98894; // @[Mux.scala 31:69:@42516.4]
  wire [15:0] _T_98895; // @[Mux.scala 31:69:@42517.4]
  wire [15:0] _T_98896; // @[Mux.scala 31:69:@42518.4]
  wire [15:0] _T_98897; // @[Mux.scala 31:69:@42519.4]
  wire [15:0] _T_98898; // @[Mux.scala 31:69:@42520.4]
  wire [15:0] _T_98899; // @[Mux.scala 31:69:@42521.4]
  wire [15:0] _T_98900; // @[Mux.scala 31:69:@42522.4]
  wire [15:0] _T_98901; // @[Mux.scala 31:69:@42523.4]
  wire  _T_98902; // @[OneHot.scala 66:30:@42524.4]
  wire  _T_98903; // @[OneHot.scala 66:30:@42525.4]
  wire  _T_98904; // @[OneHot.scala 66:30:@42526.4]
  wire  _T_98905; // @[OneHot.scala 66:30:@42527.4]
  wire  _T_98906; // @[OneHot.scala 66:30:@42528.4]
  wire  _T_98907; // @[OneHot.scala 66:30:@42529.4]
  wire  _T_98908; // @[OneHot.scala 66:30:@42530.4]
  wire  _T_98909; // @[OneHot.scala 66:30:@42531.4]
  wire  _T_98910; // @[OneHot.scala 66:30:@42532.4]
  wire  _T_98911; // @[OneHot.scala 66:30:@42533.4]
  wire  _T_98912; // @[OneHot.scala 66:30:@42534.4]
  wire  _T_98913; // @[OneHot.scala 66:30:@42535.4]
  wire  _T_98914; // @[OneHot.scala 66:30:@42536.4]
  wire  _T_98915; // @[OneHot.scala 66:30:@42537.4]
  wire  _T_98916; // @[OneHot.scala 66:30:@42538.4]
  wire  _T_98917; // @[OneHot.scala 66:30:@42539.4]
  wire [15:0] _T_98958; // @[Mux.scala 31:69:@42557.4]
  wire [15:0] _T_98959; // @[Mux.scala 31:69:@42558.4]
  wire [15:0] _T_98960; // @[Mux.scala 31:69:@42559.4]
  wire [15:0] _T_98961; // @[Mux.scala 31:69:@42560.4]
  wire [15:0] _T_98962; // @[Mux.scala 31:69:@42561.4]
  wire [15:0] _T_98963; // @[Mux.scala 31:69:@42562.4]
  wire [15:0] _T_98964; // @[Mux.scala 31:69:@42563.4]
  wire [15:0] _T_98965; // @[Mux.scala 31:69:@42564.4]
  wire [15:0] _T_98966; // @[Mux.scala 31:69:@42565.4]
  wire [15:0] _T_98967; // @[Mux.scala 31:69:@42566.4]
  wire [15:0] _T_98968; // @[Mux.scala 31:69:@42567.4]
  wire [15:0] _T_98969; // @[Mux.scala 31:69:@42568.4]
  wire [15:0] _T_98970; // @[Mux.scala 31:69:@42569.4]
  wire [15:0] _T_98971; // @[Mux.scala 31:69:@42570.4]
  wire [15:0] _T_98972; // @[Mux.scala 31:69:@42571.4]
  wire [15:0] _T_98973; // @[Mux.scala 31:69:@42572.4]
  wire  _T_98974; // @[OneHot.scala 66:30:@42573.4]
  wire  _T_98975; // @[OneHot.scala 66:30:@42574.4]
  wire  _T_98976; // @[OneHot.scala 66:30:@42575.4]
  wire  _T_98977; // @[OneHot.scala 66:30:@42576.4]
  wire  _T_98978; // @[OneHot.scala 66:30:@42577.4]
  wire  _T_98979; // @[OneHot.scala 66:30:@42578.4]
  wire  _T_98980; // @[OneHot.scala 66:30:@42579.4]
  wire  _T_98981; // @[OneHot.scala 66:30:@42580.4]
  wire  _T_98982; // @[OneHot.scala 66:30:@42581.4]
  wire  _T_98983; // @[OneHot.scala 66:30:@42582.4]
  wire  _T_98984; // @[OneHot.scala 66:30:@42583.4]
  wire  _T_98985; // @[OneHot.scala 66:30:@42584.4]
  wire  _T_98986; // @[OneHot.scala 66:30:@42585.4]
  wire  _T_98987; // @[OneHot.scala 66:30:@42586.4]
  wire  _T_98988; // @[OneHot.scala 66:30:@42587.4]
  wire  _T_98989; // @[OneHot.scala 66:30:@42588.4]
  wire [15:0] _T_99030; // @[Mux.scala 31:69:@42606.4]
  wire [15:0] _T_99031; // @[Mux.scala 31:69:@42607.4]
  wire [15:0] _T_99032; // @[Mux.scala 31:69:@42608.4]
  wire [15:0] _T_99033; // @[Mux.scala 31:69:@42609.4]
  wire [15:0] _T_99034; // @[Mux.scala 31:69:@42610.4]
  wire [15:0] _T_99035; // @[Mux.scala 31:69:@42611.4]
  wire [15:0] _T_99036; // @[Mux.scala 31:69:@42612.4]
  wire [15:0] _T_99037; // @[Mux.scala 31:69:@42613.4]
  wire [15:0] _T_99038; // @[Mux.scala 31:69:@42614.4]
  wire [15:0] _T_99039; // @[Mux.scala 31:69:@42615.4]
  wire [15:0] _T_99040; // @[Mux.scala 31:69:@42616.4]
  wire [15:0] _T_99041; // @[Mux.scala 31:69:@42617.4]
  wire [15:0] _T_99042; // @[Mux.scala 31:69:@42618.4]
  wire [15:0] _T_99043; // @[Mux.scala 31:69:@42619.4]
  wire [15:0] _T_99044; // @[Mux.scala 31:69:@42620.4]
  wire [15:0] _T_99045; // @[Mux.scala 31:69:@42621.4]
  wire  _T_99046; // @[OneHot.scala 66:30:@42622.4]
  wire  _T_99047; // @[OneHot.scala 66:30:@42623.4]
  wire  _T_99048; // @[OneHot.scala 66:30:@42624.4]
  wire  _T_99049; // @[OneHot.scala 66:30:@42625.4]
  wire  _T_99050; // @[OneHot.scala 66:30:@42626.4]
  wire  _T_99051; // @[OneHot.scala 66:30:@42627.4]
  wire  _T_99052; // @[OneHot.scala 66:30:@42628.4]
  wire  _T_99053; // @[OneHot.scala 66:30:@42629.4]
  wire  _T_99054; // @[OneHot.scala 66:30:@42630.4]
  wire  _T_99055; // @[OneHot.scala 66:30:@42631.4]
  wire  _T_99056; // @[OneHot.scala 66:30:@42632.4]
  wire  _T_99057; // @[OneHot.scala 66:30:@42633.4]
  wire  _T_99058; // @[OneHot.scala 66:30:@42634.4]
  wire  _T_99059; // @[OneHot.scala 66:30:@42635.4]
  wire  _T_99060; // @[OneHot.scala 66:30:@42636.4]
  wire  _T_99061; // @[OneHot.scala 66:30:@42637.4]
  wire [7:0] _T_99126; // @[Mux.scala 19:72:@42661.4]
  wire [15:0] _T_99134; // @[Mux.scala 19:72:@42669.4]
  wire [15:0] _T_99136; // @[Mux.scala 19:72:@42670.4]
  wire [7:0] _T_99143; // @[Mux.scala 19:72:@42677.4]
  wire [15:0] _T_99151; // @[Mux.scala 19:72:@42685.4]
  wire [15:0] _T_99153; // @[Mux.scala 19:72:@42686.4]
  wire [7:0] _T_99160; // @[Mux.scala 19:72:@42693.4]
  wire [15:0] _T_99168; // @[Mux.scala 19:72:@42701.4]
  wire [15:0] _T_99170; // @[Mux.scala 19:72:@42702.4]
  wire [7:0] _T_99177; // @[Mux.scala 19:72:@42709.4]
  wire [15:0] _T_99185; // @[Mux.scala 19:72:@42717.4]
  wire [15:0] _T_99187; // @[Mux.scala 19:72:@42718.4]
  wire [7:0] _T_99194; // @[Mux.scala 19:72:@42725.4]
  wire [15:0] _T_99202; // @[Mux.scala 19:72:@42733.4]
  wire [15:0] _T_99204; // @[Mux.scala 19:72:@42734.4]
  wire [7:0] _T_99211; // @[Mux.scala 19:72:@42741.4]
  wire [15:0] _T_99219; // @[Mux.scala 19:72:@42749.4]
  wire [15:0] _T_99221; // @[Mux.scala 19:72:@42750.4]
  wire [7:0] _T_99228; // @[Mux.scala 19:72:@42757.4]
  wire [15:0] _T_99236; // @[Mux.scala 19:72:@42765.4]
  wire [15:0] _T_99238; // @[Mux.scala 19:72:@42766.4]
  wire [7:0] _T_99245; // @[Mux.scala 19:72:@42773.4]
  wire [15:0] _T_99253; // @[Mux.scala 19:72:@42781.4]
  wire [15:0] _T_99255; // @[Mux.scala 19:72:@42782.4]
  wire [7:0] _T_99262; // @[Mux.scala 19:72:@42789.4]
  wire [15:0] _T_99270; // @[Mux.scala 19:72:@42797.4]
  wire [15:0] _T_99272; // @[Mux.scala 19:72:@42798.4]
  wire [7:0] _T_99279; // @[Mux.scala 19:72:@42805.4]
  wire [15:0] _T_99287; // @[Mux.scala 19:72:@42813.4]
  wire [15:0] _T_99289; // @[Mux.scala 19:72:@42814.4]
  wire [7:0] _T_99296; // @[Mux.scala 19:72:@42821.4]
  wire [15:0] _T_99304; // @[Mux.scala 19:72:@42829.4]
  wire [15:0] _T_99306; // @[Mux.scala 19:72:@42830.4]
  wire [7:0] _T_99313; // @[Mux.scala 19:72:@42837.4]
  wire [15:0] _T_99321; // @[Mux.scala 19:72:@42845.4]
  wire [15:0] _T_99323; // @[Mux.scala 19:72:@42846.4]
  wire [7:0] _T_99330; // @[Mux.scala 19:72:@42853.4]
  wire [15:0] _T_99338; // @[Mux.scala 19:72:@42861.4]
  wire [15:0] _T_99340; // @[Mux.scala 19:72:@42862.4]
  wire [7:0] _T_99347; // @[Mux.scala 19:72:@42869.4]
  wire [15:0] _T_99355; // @[Mux.scala 19:72:@42877.4]
  wire [15:0] _T_99357; // @[Mux.scala 19:72:@42878.4]
  wire [7:0] _T_99364; // @[Mux.scala 19:72:@42885.4]
  wire [15:0] _T_99372; // @[Mux.scala 19:72:@42893.4]
  wire [15:0] _T_99374; // @[Mux.scala 19:72:@42894.4]
  wire [7:0] _T_99381; // @[Mux.scala 19:72:@42901.4]
  wire [15:0] _T_99389; // @[Mux.scala 19:72:@42909.4]
  wire [15:0] _T_99391; // @[Mux.scala 19:72:@42910.4]
  wire [15:0] _T_99392; // @[Mux.scala 19:72:@42911.4]
  wire [15:0] _T_99393; // @[Mux.scala 19:72:@42912.4]
  wire [15:0] _T_99394; // @[Mux.scala 19:72:@42913.4]
  wire [15:0] _T_99395; // @[Mux.scala 19:72:@42914.4]
  wire [15:0] _T_99396; // @[Mux.scala 19:72:@42915.4]
  wire [15:0] _T_99397; // @[Mux.scala 19:72:@42916.4]
  wire [15:0] _T_99398; // @[Mux.scala 19:72:@42917.4]
  wire [15:0] _T_99399; // @[Mux.scala 19:72:@42918.4]
  wire [15:0] _T_99400; // @[Mux.scala 19:72:@42919.4]
  wire [15:0] _T_99401; // @[Mux.scala 19:72:@42920.4]
  wire [15:0] _T_99402; // @[Mux.scala 19:72:@42921.4]
  wire [15:0] _T_99403; // @[Mux.scala 19:72:@42922.4]
  wire [15:0] _T_99404; // @[Mux.scala 19:72:@42923.4]
  wire [15:0] _T_99405; // @[Mux.scala 19:72:@42924.4]
  wire [15:0] _T_99406; // @[Mux.scala 19:72:@42925.4]
  wire  inputPriorityPorts_1_0; // @[Mux.scala 19:72:@42929.4]
  wire  inputPriorityPorts_1_1; // @[Mux.scala 19:72:@42931.4]
  wire  inputPriorityPorts_1_2; // @[Mux.scala 19:72:@42933.4]
  wire  inputPriorityPorts_1_3; // @[Mux.scala 19:72:@42935.4]
  wire  inputPriorityPorts_1_4; // @[Mux.scala 19:72:@42937.4]
  wire  inputPriorityPorts_1_5; // @[Mux.scala 19:72:@42939.4]
  wire  inputPriorityPorts_1_6; // @[Mux.scala 19:72:@42941.4]
  wire  inputPriorityPorts_1_7; // @[Mux.scala 19:72:@42943.4]
  wire  inputPriorityPorts_1_8; // @[Mux.scala 19:72:@42945.4]
  wire  inputPriorityPorts_1_9; // @[Mux.scala 19:72:@42947.4]
  wire  inputPriorityPorts_1_10; // @[Mux.scala 19:72:@42949.4]
  wire  inputPriorityPorts_1_11; // @[Mux.scala 19:72:@42951.4]
  wire  inputPriorityPorts_1_12; // @[Mux.scala 19:72:@42953.4]
  wire  inputPriorityPorts_1_13; // @[Mux.scala 19:72:@42955.4]
  wire  inputPriorityPorts_1_14; // @[Mux.scala 19:72:@42957.4]
  wire  inputPriorityPorts_1_15; // @[Mux.scala 19:72:@42959.4]
  wire [15:0] _T_99608; // @[Mux.scala 31:69:@43013.4]
  wire [15:0] _T_99609; // @[Mux.scala 31:69:@43014.4]
  wire [15:0] _T_99610; // @[Mux.scala 31:69:@43015.4]
  wire [15:0] _T_99611; // @[Mux.scala 31:69:@43016.4]
  wire [15:0] _T_99612; // @[Mux.scala 31:69:@43017.4]
  wire [15:0] _T_99613; // @[Mux.scala 31:69:@43018.4]
  wire [15:0] _T_99614; // @[Mux.scala 31:69:@43019.4]
  wire [15:0] _T_99615; // @[Mux.scala 31:69:@43020.4]
  wire [15:0] _T_99616; // @[Mux.scala 31:69:@43021.4]
  wire [15:0] _T_99617; // @[Mux.scala 31:69:@43022.4]
  wire [15:0] _T_99618; // @[Mux.scala 31:69:@43023.4]
  wire [15:0] _T_99619; // @[Mux.scala 31:69:@43024.4]
  wire [15:0] _T_99620; // @[Mux.scala 31:69:@43025.4]
  wire [15:0] _T_99621; // @[Mux.scala 31:69:@43026.4]
  wire [15:0] _T_99622; // @[Mux.scala 31:69:@43027.4]
  wire [15:0] _T_99623; // @[Mux.scala 31:69:@43028.4]
  wire  _T_99624; // @[OneHot.scala 66:30:@43029.4]
  wire  _T_99625; // @[OneHot.scala 66:30:@43030.4]
  wire  _T_99626; // @[OneHot.scala 66:30:@43031.4]
  wire  _T_99627; // @[OneHot.scala 66:30:@43032.4]
  wire  _T_99628; // @[OneHot.scala 66:30:@43033.4]
  wire  _T_99629; // @[OneHot.scala 66:30:@43034.4]
  wire  _T_99630; // @[OneHot.scala 66:30:@43035.4]
  wire  _T_99631; // @[OneHot.scala 66:30:@43036.4]
  wire  _T_99632; // @[OneHot.scala 66:30:@43037.4]
  wire  _T_99633; // @[OneHot.scala 66:30:@43038.4]
  wire  _T_99634; // @[OneHot.scala 66:30:@43039.4]
  wire  _T_99635; // @[OneHot.scala 66:30:@43040.4]
  wire  _T_99636; // @[OneHot.scala 66:30:@43041.4]
  wire  _T_99637; // @[OneHot.scala 66:30:@43042.4]
  wire  _T_99638; // @[OneHot.scala 66:30:@43043.4]
  wire  _T_99639; // @[OneHot.scala 66:30:@43044.4]
  wire [15:0] _T_99680; // @[Mux.scala 31:69:@43062.4]
  wire [15:0] _T_99681; // @[Mux.scala 31:69:@43063.4]
  wire [15:0] _T_99682; // @[Mux.scala 31:69:@43064.4]
  wire [15:0] _T_99683; // @[Mux.scala 31:69:@43065.4]
  wire [15:0] _T_99684; // @[Mux.scala 31:69:@43066.4]
  wire [15:0] _T_99685; // @[Mux.scala 31:69:@43067.4]
  wire [15:0] _T_99686; // @[Mux.scala 31:69:@43068.4]
  wire [15:0] _T_99687; // @[Mux.scala 31:69:@43069.4]
  wire [15:0] _T_99688; // @[Mux.scala 31:69:@43070.4]
  wire [15:0] _T_99689; // @[Mux.scala 31:69:@43071.4]
  wire [15:0] _T_99690; // @[Mux.scala 31:69:@43072.4]
  wire [15:0] _T_99691; // @[Mux.scala 31:69:@43073.4]
  wire [15:0] _T_99692; // @[Mux.scala 31:69:@43074.4]
  wire [15:0] _T_99693; // @[Mux.scala 31:69:@43075.4]
  wire [15:0] _T_99694; // @[Mux.scala 31:69:@43076.4]
  wire [15:0] _T_99695; // @[Mux.scala 31:69:@43077.4]
  wire  _T_99696; // @[OneHot.scala 66:30:@43078.4]
  wire  _T_99697; // @[OneHot.scala 66:30:@43079.4]
  wire  _T_99698; // @[OneHot.scala 66:30:@43080.4]
  wire  _T_99699; // @[OneHot.scala 66:30:@43081.4]
  wire  _T_99700; // @[OneHot.scala 66:30:@43082.4]
  wire  _T_99701; // @[OneHot.scala 66:30:@43083.4]
  wire  _T_99702; // @[OneHot.scala 66:30:@43084.4]
  wire  _T_99703; // @[OneHot.scala 66:30:@43085.4]
  wire  _T_99704; // @[OneHot.scala 66:30:@43086.4]
  wire  _T_99705; // @[OneHot.scala 66:30:@43087.4]
  wire  _T_99706; // @[OneHot.scala 66:30:@43088.4]
  wire  _T_99707; // @[OneHot.scala 66:30:@43089.4]
  wire  _T_99708; // @[OneHot.scala 66:30:@43090.4]
  wire  _T_99709; // @[OneHot.scala 66:30:@43091.4]
  wire  _T_99710; // @[OneHot.scala 66:30:@43092.4]
  wire  _T_99711; // @[OneHot.scala 66:30:@43093.4]
  wire [15:0] _T_99752; // @[Mux.scala 31:69:@43111.4]
  wire [15:0] _T_99753; // @[Mux.scala 31:69:@43112.4]
  wire [15:0] _T_99754; // @[Mux.scala 31:69:@43113.4]
  wire [15:0] _T_99755; // @[Mux.scala 31:69:@43114.4]
  wire [15:0] _T_99756; // @[Mux.scala 31:69:@43115.4]
  wire [15:0] _T_99757; // @[Mux.scala 31:69:@43116.4]
  wire [15:0] _T_99758; // @[Mux.scala 31:69:@43117.4]
  wire [15:0] _T_99759; // @[Mux.scala 31:69:@43118.4]
  wire [15:0] _T_99760; // @[Mux.scala 31:69:@43119.4]
  wire [15:0] _T_99761; // @[Mux.scala 31:69:@43120.4]
  wire [15:0] _T_99762; // @[Mux.scala 31:69:@43121.4]
  wire [15:0] _T_99763; // @[Mux.scala 31:69:@43122.4]
  wire [15:0] _T_99764; // @[Mux.scala 31:69:@43123.4]
  wire [15:0] _T_99765; // @[Mux.scala 31:69:@43124.4]
  wire [15:0] _T_99766; // @[Mux.scala 31:69:@43125.4]
  wire [15:0] _T_99767; // @[Mux.scala 31:69:@43126.4]
  wire  _T_99768; // @[OneHot.scala 66:30:@43127.4]
  wire  _T_99769; // @[OneHot.scala 66:30:@43128.4]
  wire  _T_99770; // @[OneHot.scala 66:30:@43129.4]
  wire  _T_99771; // @[OneHot.scala 66:30:@43130.4]
  wire  _T_99772; // @[OneHot.scala 66:30:@43131.4]
  wire  _T_99773; // @[OneHot.scala 66:30:@43132.4]
  wire  _T_99774; // @[OneHot.scala 66:30:@43133.4]
  wire  _T_99775; // @[OneHot.scala 66:30:@43134.4]
  wire  _T_99776; // @[OneHot.scala 66:30:@43135.4]
  wire  _T_99777; // @[OneHot.scala 66:30:@43136.4]
  wire  _T_99778; // @[OneHot.scala 66:30:@43137.4]
  wire  _T_99779; // @[OneHot.scala 66:30:@43138.4]
  wire  _T_99780; // @[OneHot.scala 66:30:@43139.4]
  wire  _T_99781; // @[OneHot.scala 66:30:@43140.4]
  wire  _T_99782; // @[OneHot.scala 66:30:@43141.4]
  wire  _T_99783; // @[OneHot.scala 66:30:@43142.4]
  wire [15:0] _T_99824; // @[Mux.scala 31:69:@43160.4]
  wire [15:0] _T_99825; // @[Mux.scala 31:69:@43161.4]
  wire [15:0] _T_99826; // @[Mux.scala 31:69:@43162.4]
  wire [15:0] _T_99827; // @[Mux.scala 31:69:@43163.4]
  wire [15:0] _T_99828; // @[Mux.scala 31:69:@43164.4]
  wire [15:0] _T_99829; // @[Mux.scala 31:69:@43165.4]
  wire [15:0] _T_99830; // @[Mux.scala 31:69:@43166.4]
  wire [15:0] _T_99831; // @[Mux.scala 31:69:@43167.4]
  wire [15:0] _T_99832; // @[Mux.scala 31:69:@43168.4]
  wire [15:0] _T_99833; // @[Mux.scala 31:69:@43169.4]
  wire [15:0] _T_99834; // @[Mux.scala 31:69:@43170.4]
  wire [15:0] _T_99835; // @[Mux.scala 31:69:@43171.4]
  wire [15:0] _T_99836; // @[Mux.scala 31:69:@43172.4]
  wire [15:0] _T_99837; // @[Mux.scala 31:69:@43173.4]
  wire [15:0] _T_99838; // @[Mux.scala 31:69:@43174.4]
  wire [15:0] _T_99839; // @[Mux.scala 31:69:@43175.4]
  wire  _T_99840; // @[OneHot.scala 66:30:@43176.4]
  wire  _T_99841; // @[OneHot.scala 66:30:@43177.4]
  wire  _T_99842; // @[OneHot.scala 66:30:@43178.4]
  wire  _T_99843; // @[OneHot.scala 66:30:@43179.4]
  wire  _T_99844; // @[OneHot.scala 66:30:@43180.4]
  wire  _T_99845; // @[OneHot.scala 66:30:@43181.4]
  wire  _T_99846; // @[OneHot.scala 66:30:@43182.4]
  wire  _T_99847; // @[OneHot.scala 66:30:@43183.4]
  wire  _T_99848; // @[OneHot.scala 66:30:@43184.4]
  wire  _T_99849; // @[OneHot.scala 66:30:@43185.4]
  wire  _T_99850; // @[OneHot.scala 66:30:@43186.4]
  wire  _T_99851; // @[OneHot.scala 66:30:@43187.4]
  wire  _T_99852; // @[OneHot.scala 66:30:@43188.4]
  wire  _T_99853; // @[OneHot.scala 66:30:@43189.4]
  wire  _T_99854; // @[OneHot.scala 66:30:@43190.4]
  wire  _T_99855; // @[OneHot.scala 66:30:@43191.4]
  wire [15:0] _T_99896; // @[Mux.scala 31:69:@43209.4]
  wire [15:0] _T_99897; // @[Mux.scala 31:69:@43210.4]
  wire [15:0] _T_99898; // @[Mux.scala 31:69:@43211.4]
  wire [15:0] _T_99899; // @[Mux.scala 31:69:@43212.4]
  wire [15:0] _T_99900; // @[Mux.scala 31:69:@43213.4]
  wire [15:0] _T_99901; // @[Mux.scala 31:69:@43214.4]
  wire [15:0] _T_99902; // @[Mux.scala 31:69:@43215.4]
  wire [15:0] _T_99903; // @[Mux.scala 31:69:@43216.4]
  wire [15:0] _T_99904; // @[Mux.scala 31:69:@43217.4]
  wire [15:0] _T_99905; // @[Mux.scala 31:69:@43218.4]
  wire [15:0] _T_99906; // @[Mux.scala 31:69:@43219.4]
  wire [15:0] _T_99907; // @[Mux.scala 31:69:@43220.4]
  wire [15:0] _T_99908; // @[Mux.scala 31:69:@43221.4]
  wire [15:0] _T_99909; // @[Mux.scala 31:69:@43222.4]
  wire [15:0] _T_99910; // @[Mux.scala 31:69:@43223.4]
  wire [15:0] _T_99911; // @[Mux.scala 31:69:@43224.4]
  wire  _T_99912; // @[OneHot.scala 66:30:@43225.4]
  wire  _T_99913; // @[OneHot.scala 66:30:@43226.4]
  wire  _T_99914; // @[OneHot.scala 66:30:@43227.4]
  wire  _T_99915; // @[OneHot.scala 66:30:@43228.4]
  wire  _T_99916; // @[OneHot.scala 66:30:@43229.4]
  wire  _T_99917; // @[OneHot.scala 66:30:@43230.4]
  wire  _T_99918; // @[OneHot.scala 66:30:@43231.4]
  wire  _T_99919; // @[OneHot.scala 66:30:@43232.4]
  wire  _T_99920; // @[OneHot.scala 66:30:@43233.4]
  wire  _T_99921; // @[OneHot.scala 66:30:@43234.4]
  wire  _T_99922; // @[OneHot.scala 66:30:@43235.4]
  wire  _T_99923; // @[OneHot.scala 66:30:@43236.4]
  wire  _T_99924; // @[OneHot.scala 66:30:@43237.4]
  wire  _T_99925; // @[OneHot.scala 66:30:@43238.4]
  wire  _T_99926; // @[OneHot.scala 66:30:@43239.4]
  wire  _T_99927; // @[OneHot.scala 66:30:@43240.4]
  wire [15:0] _T_99968; // @[Mux.scala 31:69:@43258.4]
  wire [15:0] _T_99969; // @[Mux.scala 31:69:@43259.4]
  wire [15:0] _T_99970; // @[Mux.scala 31:69:@43260.4]
  wire [15:0] _T_99971; // @[Mux.scala 31:69:@43261.4]
  wire [15:0] _T_99972; // @[Mux.scala 31:69:@43262.4]
  wire [15:0] _T_99973; // @[Mux.scala 31:69:@43263.4]
  wire [15:0] _T_99974; // @[Mux.scala 31:69:@43264.4]
  wire [15:0] _T_99975; // @[Mux.scala 31:69:@43265.4]
  wire [15:0] _T_99976; // @[Mux.scala 31:69:@43266.4]
  wire [15:0] _T_99977; // @[Mux.scala 31:69:@43267.4]
  wire [15:0] _T_99978; // @[Mux.scala 31:69:@43268.4]
  wire [15:0] _T_99979; // @[Mux.scala 31:69:@43269.4]
  wire [15:0] _T_99980; // @[Mux.scala 31:69:@43270.4]
  wire [15:0] _T_99981; // @[Mux.scala 31:69:@43271.4]
  wire [15:0] _T_99982; // @[Mux.scala 31:69:@43272.4]
  wire [15:0] _T_99983; // @[Mux.scala 31:69:@43273.4]
  wire  _T_99984; // @[OneHot.scala 66:30:@43274.4]
  wire  _T_99985; // @[OneHot.scala 66:30:@43275.4]
  wire  _T_99986; // @[OneHot.scala 66:30:@43276.4]
  wire  _T_99987; // @[OneHot.scala 66:30:@43277.4]
  wire  _T_99988; // @[OneHot.scala 66:30:@43278.4]
  wire  _T_99989; // @[OneHot.scala 66:30:@43279.4]
  wire  _T_99990; // @[OneHot.scala 66:30:@43280.4]
  wire  _T_99991; // @[OneHot.scala 66:30:@43281.4]
  wire  _T_99992; // @[OneHot.scala 66:30:@43282.4]
  wire  _T_99993; // @[OneHot.scala 66:30:@43283.4]
  wire  _T_99994; // @[OneHot.scala 66:30:@43284.4]
  wire  _T_99995; // @[OneHot.scala 66:30:@43285.4]
  wire  _T_99996; // @[OneHot.scala 66:30:@43286.4]
  wire  _T_99997; // @[OneHot.scala 66:30:@43287.4]
  wire  _T_99998; // @[OneHot.scala 66:30:@43288.4]
  wire  _T_99999; // @[OneHot.scala 66:30:@43289.4]
  wire [15:0] _T_100040; // @[Mux.scala 31:69:@43307.4]
  wire [15:0] _T_100041; // @[Mux.scala 31:69:@43308.4]
  wire [15:0] _T_100042; // @[Mux.scala 31:69:@43309.4]
  wire [15:0] _T_100043; // @[Mux.scala 31:69:@43310.4]
  wire [15:0] _T_100044; // @[Mux.scala 31:69:@43311.4]
  wire [15:0] _T_100045; // @[Mux.scala 31:69:@43312.4]
  wire [15:0] _T_100046; // @[Mux.scala 31:69:@43313.4]
  wire [15:0] _T_100047; // @[Mux.scala 31:69:@43314.4]
  wire [15:0] _T_100048; // @[Mux.scala 31:69:@43315.4]
  wire [15:0] _T_100049; // @[Mux.scala 31:69:@43316.4]
  wire [15:0] _T_100050; // @[Mux.scala 31:69:@43317.4]
  wire [15:0] _T_100051; // @[Mux.scala 31:69:@43318.4]
  wire [15:0] _T_100052; // @[Mux.scala 31:69:@43319.4]
  wire [15:0] _T_100053; // @[Mux.scala 31:69:@43320.4]
  wire [15:0] _T_100054; // @[Mux.scala 31:69:@43321.4]
  wire [15:0] _T_100055; // @[Mux.scala 31:69:@43322.4]
  wire  _T_100056; // @[OneHot.scala 66:30:@43323.4]
  wire  _T_100057; // @[OneHot.scala 66:30:@43324.4]
  wire  _T_100058; // @[OneHot.scala 66:30:@43325.4]
  wire  _T_100059; // @[OneHot.scala 66:30:@43326.4]
  wire  _T_100060; // @[OneHot.scala 66:30:@43327.4]
  wire  _T_100061; // @[OneHot.scala 66:30:@43328.4]
  wire  _T_100062; // @[OneHot.scala 66:30:@43329.4]
  wire  _T_100063; // @[OneHot.scala 66:30:@43330.4]
  wire  _T_100064; // @[OneHot.scala 66:30:@43331.4]
  wire  _T_100065; // @[OneHot.scala 66:30:@43332.4]
  wire  _T_100066; // @[OneHot.scala 66:30:@43333.4]
  wire  _T_100067; // @[OneHot.scala 66:30:@43334.4]
  wire  _T_100068; // @[OneHot.scala 66:30:@43335.4]
  wire  _T_100069; // @[OneHot.scala 66:30:@43336.4]
  wire  _T_100070; // @[OneHot.scala 66:30:@43337.4]
  wire  _T_100071; // @[OneHot.scala 66:30:@43338.4]
  wire [15:0] _T_100112; // @[Mux.scala 31:69:@43356.4]
  wire [15:0] _T_100113; // @[Mux.scala 31:69:@43357.4]
  wire [15:0] _T_100114; // @[Mux.scala 31:69:@43358.4]
  wire [15:0] _T_100115; // @[Mux.scala 31:69:@43359.4]
  wire [15:0] _T_100116; // @[Mux.scala 31:69:@43360.4]
  wire [15:0] _T_100117; // @[Mux.scala 31:69:@43361.4]
  wire [15:0] _T_100118; // @[Mux.scala 31:69:@43362.4]
  wire [15:0] _T_100119; // @[Mux.scala 31:69:@43363.4]
  wire [15:0] _T_100120; // @[Mux.scala 31:69:@43364.4]
  wire [15:0] _T_100121; // @[Mux.scala 31:69:@43365.4]
  wire [15:0] _T_100122; // @[Mux.scala 31:69:@43366.4]
  wire [15:0] _T_100123; // @[Mux.scala 31:69:@43367.4]
  wire [15:0] _T_100124; // @[Mux.scala 31:69:@43368.4]
  wire [15:0] _T_100125; // @[Mux.scala 31:69:@43369.4]
  wire [15:0] _T_100126; // @[Mux.scala 31:69:@43370.4]
  wire [15:0] _T_100127; // @[Mux.scala 31:69:@43371.4]
  wire  _T_100128; // @[OneHot.scala 66:30:@43372.4]
  wire  _T_100129; // @[OneHot.scala 66:30:@43373.4]
  wire  _T_100130; // @[OneHot.scala 66:30:@43374.4]
  wire  _T_100131; // @[OneHot.scala 66:30:@43375.4]
  wire  _T_100132; // @[OneHot.scala 66:30:@43376.4]
  wire  _T_100133; // @[OneHot.scala 66:30:@43377.4]
  wire  _T_100134; // @[OneHot.scala 66:30:@43378.4]
  wire  _T_100135; // @[OneHot.scala 66:30:@43379.4]
  wire  _T_100136; // @[OneHot.scala 66:30:@43380.4]
  wire  _T_100137; // @[OneHot.scala 66:30:@43381.4]
  wire  _T_100138; // @[OneHot.scala 66:30:@43382.4]
  wire  _T_100139; // @[OneHot.scala 66:30:@43383.4]
  wire  _T_100140; // @[OneHot.scala 66:30:@43384.4]
  wire  _T_100141; // @[OneHot.scala 66:30:@43385.4]
  wire  _T_100142; // @[OneHot.scala 66:30:@43386.4]
  wire  _T_100143; // @[OneHot.scala 66:30:@43387.4]
  wire [15:0] _T_100184; // @[Mux.scala 31:69:@43405.4]
  wire [15:0] _T_100185; // @[Mux.scala 31:69:@43406.4]
  wire [15:0] _T_100186; // @[Mux.scala 31:69:@43407.4]
  wire [15:0] _T_100187; // @[Mux.scala 31:69:@43408.4]
  wire [15:0] _T_100188; // @[Mux.scala 31:69:@43409.4]
  wire [15:0] _T_100189; // @[Mux.scala 31:69:@43410.4]
  wire [15:0] _T_100190; // @[Mux.scala 31:69:@43411.4]
  wire [15:0] _T_100191; // @[Mux.scala 31:69:@43412.4]
  wire [15:0] _T_100192; // @[Mux.scala 31:69:@43413.4]
  wire [15:0] _T_100193; // @[Mux.scala 31:69:@43414.4]
  wire [15:0] _T_100194; // @[Mux.scala 31:69:@43415.4]
  wire [15:0] _T_100195; // @[Mux.scala 31:69:@43416.4]
  wire [15:0] _T_100196; // @[Mux.scala 31:69:@43417.4]
  wire [15:0] _T_100197; // @[Mux.scala 31:69:@43418.4]
  wire [15:0] _T_100198; // @[Mux.scala 31:69:@43419.4]
  wire [15:0] _T_100199; // @[Mux.scala 31:69:@43420.4]
  wire  _T_100200; // @[OneHot.scala 66:30:@43421.4]
  wire  _T_100201; // @[OneHot.scala 66:30:@43422.4]
  wire  _T_100202; // @[OneHot.scala 66:30:@43423.4]
  wire  _T_100203; // @[OneHot.scala 66:30:@43424.4]
  wire  _T_100204; // @[OneHot.scala 66:30:@43425.4]
  wire  _T_100205; // @[OneHot.scala 66:30:@43426.4]
  wire  _T_100206; // @[OneHot.scala 66:30:@43427.4]
  wire  _T_100207; // @[OneHot.scala 66:30:@43428.4]
  wire  _T_100208; // @[OneHot.scala 66:30:@43429.4]
  wire  _T_100209; // @[OneHot.scala 66:30:@43430.4]
  wire  _T_100210; // @[OneHot.scala 66:30:@43431.4]
  wire  _T_100211; // @[OneHot.scala 66:30:@43432.4]
  wire  _T_100212; // @[OneHot.scala 66:30:@43433.4]
  wire  _T_100213; // @[OneHot.scala 66:30:@43434.4]
  wire  _T_100214; // @[OneHot.scala 66:30:@43435.4]
  wire  _T_100215; // @[OneHot.scala 66:30:@43436.4]
  wire [15:0] _T_100256; // @[Mux.scala 31:69:@43454.4]
  wire [15:0] _T_100257; // @[Mux.scala 31:69:@43455.4]
  wire [15:0] _T_100258; // @[Mux.scala 31:69:@43456.4]
  wire [15:0] _T_100259; // @[Mux.scala 31:69:@43457.4]
  wire [15:0] _T_100260; // @[Mux.scala 31:69:@43458.4]
  wire [15:0] _T_100261; // @[Mux.scala 31:69:@43459.4]
  wire [15:0] _T_100262; // @[Mux.scala 31:69:@43460.4]
  wire [15:0] _T_100263; // @[Mux.scala 31:69:@43461.4]
  wire [15:0] _T_100264; // @[Mux.scala 31:69:@43462.4]
  wire [15:0] _T_100265; // @[Mux.scala 31:69:@43463.4]
  wire [15:0] _T_100266; // @[Mux.scala 31:69:@43464.4]
  wire [15:0] _T_100267; // @[Mux.scala 31:69:@43465.4]
  wire [15:0] _T_100268; // @[Mux.scala 31:69:@43466.4]
  wire [15:0] _T_100269; // @[Mux.scala 31:69:@43467.4]
  wire [15:0] _T_100270; // @[Mux.scala 31:69:@43468.4]
  wire [15:0] _T_100271; // @[Mux.scala 31:69:@43469.4]
  wire  _T_100272; // @[OneHot.scala 66:30:@43470.4]
  wire  _T_100273; // @[OneHot.scala 66:30:@43471.4]
  wire  _T_100274; // @[OneHot.scala 66:30:@43472.4]
  wire  _T_100275; // @[OneHot.scala 66:30:@43473.4]
  wire  _T_100276; // @[OneHot.scala 66:30:@43474.4]
  wire  _T_100277; // @[OneHot.scala 66:30:@43475.4]
  wire  _T_100278; // @[OneHot.scala 66:30:@43476.4]
  wire  _T_100279; // @[OneHot.scala 66:30:@43477.4]
  wire  _T_100280; // @[OneHot.scala 66:30:@43478.4]
  wire  _T_100281; // @[OneHot.scala 66:30:@43479.4]
  wire  _T_100282; // @[OneHot.scala 66:30:@43480.4]
  wire  _T_100283; // @[OneHot.scala 66:30:@43481.4]
  wire  _T_100284; // @[OneHot.scala 66:30:@43482.4]
  wire  _T_100285; // @[OneHot.scala 66:30:@43483.4]
  wire  _T_100286; // @[OneHot.scala 66:30:@43484.4]
  wire  _T_100287; // @[OneHot.scala 66:30:@43485.4]
  wire [15:0] _T_100328; // @[Mux.scala 31:69:@43503.4]
  wire [15:0] _T_100329; // @[Mux.scala 31:69:@43504.4]
  wire [15:0] _T_100330; // @[Mux.scala 31:69:@43505.4]
  wire [15:0] _T_100331; // @[Mux.scala 31:69:@43506.4]
  wire [15:0] _T_100332; // @[Mux.scala 31:69:@43507.4]
  wire [15:0] _T_100333; // @[Mux.scala 31:69:@43508.4]
  wire [15:0] _T_100334; // @[Mux.scala 31:69:@43509.4]
  wire [15:0] _T_100335; // @[Mux.scala 31:69:@43510.4]
  wire [15:0] _T_100336; // @[Mux.scala 31:69:@43511.4]
  wire [15:0] _T_100337; // @[Mux.scala 31:69:@43512.4]
  wire [15:0] _T_100338; // @[Mux.scala 31:69:@43513.4]
  wire [15:0] _T_100339; // @[Mux.scala 31:69:@43514.4]
  wire [15:0] _T_100340; // @[Mux.scala 31:69:@43515.4]
  wire [15:0] _T_100341; // @[Mux.scala 31:69:@43516.4]
  wire [15:0] _T_100342; // @[Mux.scala 31:69:@43517.4]
  wire [15:0] _T_100343; // @[Mux.scala 31:69:@43518.4]
  wire  _T_100344; // @[OneHot.scala 66:30:@43519.4]
  wire  _T_100345; // @[OneHot.scala 66:30:@43520.4]
  wire  _T_100346; // @[OneHot.scala 66:30:@43521.4]
  wire  _T_100347; // @[OneHot.scala 66:30:@43522.4]
  wire  _T_100348; // @[OneHot.scala 66:30:@43523.4]
  wire  _T_100349; // @[OneHot.scala 66:30:@43524.4]
  wire  _T_100350; // @[OneHot.scala 66:30:@43525.4]
  wire  _T_100351; // @[OneHot.scala 66:30:@43526.4]
  wire  _T_100352; // @[OneHot.scala 66:30:@43527.4]
  wire  _T_100353; // @[OneHot.scala 66:30:@43528.4]
  wire  _T_100354; // @[OneHot.scala 66:30:@43529.4]
  wire  _T_100355; // @[OneHot.scala 66:30:@43530.4]
  wire  _T_100356; // @[OneHot.scala 66:30:@43531.4]
  wire  _T_100357; // @[OneHot.scala 66:30:@43532.4]
  wire  _T_100358; // @[OneHot.scala 66:30:@43533.4]
  wire  _T_100359; // @[OneHot.scala 66:30:@43534.4]
  wire [15:0] _T_100400; // @[Mux.scala 31:69:@43552.4]
  wire [15:0] _T_100401; // @[Mux.scala 31:69:@43553.4]
  wire [15:0] _T_100402; // @[Mux.scala 31:69:@43554.4]
  wire [15:0] _T_100403; // @[Mux.scala 31:69:@43555.4]
  wire [15:0] _T_100404; // @[Mux.scala 31:69:@43556.4]
  wire [15:0] _T_100405; // @[Mux.scala 31:69:@43557.4]
  wire [15:0] _T_100406; // @[Mux.scala 31:69:@43558.4]
  wire [15:0] _T_100407; // @[Mux.scala 31:69:@43559.4]
  wire [15:0] _T_100408; // @[Mux.scala 31:69:@43560.4]
  wire [15:0] _T_100409; // @[Mux.scala 31:69:@43561.4]
  wire [15:0] _T_100410; // @[Mux.scala 31:69:@43562.4]
  wire [15:0] _T_100411; // @[Mux.scala 31:69:@43563.4]
  wire [15:0] _T_100412; // @[Mux.scala 31:69:@43564.4]
  wire [15:0] _T_100413; // @[Mux.scala 31:69:@43565.4]
  wire [15:0] _T_100414; // @[Mux.scala 31:69:@43566.4]
  wire [15:0] _T_100415; // @[Mux.scala 31:69:@43567.4]
  wire  _T_100416; // @[OneHot.scala 66:30:@43568.4]
  wire  _T_100417; // @[OneHot.scala 66:30:@43569.4]
  wire  _T_100418; // @[OneHot.scala 66:30:@43570.4]
  wire  _T_100419; // @[OneHot.scala 66:30:@43571.4]
  wire  _T_100420; // @[OneHot.scala 66:30:@43572.4]
  wire  _T_100421; // @[OneHot.scala 66:30:@43573.4]
  wire  _T_100422; // @[OneHot.scala 66:30:@43574.4]
  wire  _T_100423; // @[OneHot.scala 66:30:@43575.4]
  wire  _T_100424; // @[OneHot.scala 66:30:@43576.4]
  wire  _T_100425; // @[OneHot.scala 66:30:@43577.4]
  wire  _T_100426; // @[OneHot.scala 66:30:@43578.4]
  wire  _T_100427; // @[OneHot.scala 66:30:@43579.4]
  wire  _T_100428; // @[OneHot.scala 66:30:@43580.4]
  wire  _T_100429; // @[OneHot.scala 66:30:@43581.4]
  wire  _T_100430; // @[OneHot.scala 66:30:@43582.4]
  wire  _T_100431; // @[OneHot.scala 66:30:@43583.4]
  wire [15:0] _T_100472; // @[Mux.scala 31:69:@43601.4]
  wire [15:0] _T_100473; // @[Mux.scala 31:69:@43602.4]
  wire [15:0] _T_100474; // @[Mux.scala 31:69:@43603.4]
  wire [15:0] _T_100475; // @[Mux.scala 31:69:@43604.4]
  wire [15:0] _T_100476; // @[Mux.scala 31:69:@43605.4]
  wire [15:0] _T_100477; // @[Mux.scala 31:69:@43606.4]
  wire [15:0] _T_100478; // @[Mux.scala 31:69:@43607.4]
  wire [15:0] _T_100479; // @[Mux.scala 31:69:@43608.4]
  wire [15:0] _T_100480; // @[Mux.scala 31:69:@43609.4]
  wire [15:0] _T_100481; // @[Mux.scala 31:69:@43610.4]
  wire [15:0] _T_100482; // @[Mux.scala 31:69:@43611.4]
  wire [15:0] _T_100483; // @[Mux.scala 31:69:@43612.4]
  wire [15:0] _T_100484; // @[Mux.scala 31:69:@43613.4]
  wire [15:0] _T_100485; // @[Mux.scala 31:69:@43614.4]
  wire [15:0] _T_100486; // @[Mux.scala 31:69:@43615.4]
  wire [15:0] _T_100487; // @[Mux.scala 31:69:@43616.4]
  wire  _T_100488; // @[OneHot.scala 66:30:@43617.4]
  wire  _T_100489; // @[OneHot.scala 66:30:@43618.4]
  wire  _T_100490; // @[OneHot.scala 66:30:@43619.4]
  wire  _T_100491; // @[OneHot.scala 66:30:@43620.4]
  wire  _T_100492; // @[OneHot.scala 66:30:@43621.4]
  wire  _T_100493; // @[OneHot.scala 66:30:@43622.4]
  wire  _T_100494; // @[OneHot.scala 66:30:@43623.4]
  wire  _T_100495; // @[OneHot.scala 66:30:@43624.4]
  wire  _T_100496; // @[OneHot.scala 66:30:@43625.4]
  wire  _T_100497; // @[OneHot.scala 66:30:@43626.4]
  wire  _T_100498; // @[OneHot.scala 66:30:@43627.4]
  wire  _T_100499; // @[OneHot.scala 66:30:@43628.4]
  wire  _T_100500; // @[OneHot.scala 66:30:@43629.4]
  wire  _T_100501; // @[OneHot.scala 66:30:@43630.4]
  wire  _T_100502; // @[OneHot.scala 66:30:@43631.4]
  wire  _T_100503; // @[OneHot.scala 66:30:@43632.4]
  wire [15:0] _T_100544; // @[Mux.scala 31:69:@43650.4]
  wire [15:0] _T_100545; // @[Mux.scala 31:69:@43651.4]
  wire [15:0] _T_100546; // @[Mux.scala 31:69:@43652.4]
  wire [15:0] _T_100547; // @[Mux.scala 31:69:@43653.4]
  wire [15:0] _T_100548; // @[Mux.scala 31:69:@43654.4]
  wire [15:0] _T_100549; // @[Mux.scala 31:69:@43655.4]
  wire [15:0] _T_100550; // @[Mux.scala 31:69:@43656.4]
  wire [15:0] _T_100551; // @[Mux.scala 31:69:@43657.4]
  wire [15:0] _T_100552; // @[Mux.scala 31:69:@43658.4]
  wire [15:0] _T_100553; // @[Mux.scala 31:69:@43659.4]
  wire [15:0] _T_100554; // @[Mux.scala 31:69:@43660.4]
  wire [15:0] _T_100555; // @[Mux.scala 31:69:@43661.4]
  wire [15:0] _T_100556; // @[Mux.scala 31:69:@43662.4]
  wire [15:0] _T_100557; // @[Mux.scala 31:69:@43663.4]
  wire [15:0] _T_100558; // @[Mux.scala 31:69:@43664.4]
  wire [15:0] _T_100559; // @[Mux.scala 31:69:@43665.4]
  wire  _T_100560; // @[OneHot.scala 66:30:@43666.4]
  wire  _T_100561; // @[OneHot.scala 66:30:@43667.4]
  wire  _T_100562; // @[OneHot.scala 66:30:@43668.4]
  wire  _T_100563; // @[OneHot.scala 66:30:@43669.4]
  wire  _T_100564; // @[OneHot.scala 66:30:@43670.4]
  wire  _T_100565; // @[OneHot.scala 66:30:@43671.4]
  wire  _T_100566; // @[OneHot.scala 66:30:@43672.4]
  wire  _T_100567; // @[OneHot.scala 66:30:@43673.4]
  wire  _T_100568; // @[OneHot.scala 66:30:@43674.4]
  wire  _T_100569; // @[OneHot.scala 66:30:@43675.4]
  wire  _T_100570; // @[OneHot.scala 66:30:@43676.4]
  wire  _T_100571; // @[OneHot.scala 66:30:@43677.4]
  wire  _T_100572; // @[OneHot.scala 66:30:@43678.4]
  wire  _T_100573; // @[OneHot.scala 66:30:@43679.4]
  wire  _T_100574; // @[OneHot.scala 66:30:@43680.4]
  wire  _T_100575; // @[OneHot.scala 66:30:@43681.4]
  wire [15:0] _T_100616; // @[Mux.scala 31:69:@43699.4]
  wire [15:0] _T_100617; // @[Mux.scala 31:69:@43700.4]
  wire [15:0] _T_100618; // @[Mux.scala 31:69:@43701.4]
  wire [15:0] _T_100619; // @[Mux.scala 31:69:@43702.4]
  wire [15:0] _T_100620; // @[Mux.scala 31:69:@43703.4]
  wire [15:0] _T_100621; // @[Mux.scala 31:69:@43704.4]
  wire [15:0] _T_100622; // @[Mux.scala 31:69:@43705.4]
  wire [15:0] _T_100623; // @[Mux.scala 31:69:@43706.4]
  wire [15:0] _T_100624; // @[Mux.scala 31:69:@43707.4]
  wire [15:0] _T_100625; // @[Mux.scala 31:69:@43708.4]
  wire [15:0] _T_100626; // @[Mux.scala 31:69:@43709.4]
  wire [15:0] _T_100627; // @[Mux.scala 31:69:@43710.4]
  wire [15:0] _T_100628; // @[Mux.scala 31:69:@43711.4]
  wire [15:0] _T_100629; // @[Mux.scala 31:69:@43712.4]
  wire [15:0] _T_100630; // @[Mux.scala 31:69:@43713.4]
  wire [15:0] _T_100631; // @[Mux.scala 31:69:@43714.4]
  wire  _T_100632; // @[OneHot.scala 66:30:@43715.4]
  wire  _T_100633; // @[OneHot.scala 66:30:@43716.4]
  wire  _T_100634; // @[OneHot.scala 66:30:@43717.4]
  wire  _T_100635; // @[OneHot.scala 66:30:@43718.4]
  wire  _T_100636; // @[OneHot.scala 66:30:@43719.4]
  wire  _T_100637; // @[OneHot.scala 66:30:@43720.4]
  wire  _T_100638; // @[OneHot.scala 66:30:@43721.4]
  wire  _T_100639; // @[OneHot.scala 66:30:@43722.4]
  wire  _T_100640; // @[OneHot.scala 66:30:@43723.4]
  wire  _T_100641; // @[OneHot.scala 66:30:@43724.4]
  wire  _T_100642; // @[OneHot.scala 66:30:@43725.4]
  wire  _T_100643; // @[OneHot.scala 66:30:@43726.4]
  wire  _T_100644; // @[OneHot.scala 66:30:@43727.4]
  wire  _T_100645; // @[OneHot.scala 66:30:@43728.4]
  wire  _T_100646; // @[OneHot.scala 66:30:@43729.4]
  wire  _T_100647; // @[OneHot.scala 66:30:@43730.4]
  wire [15:0] _T_100688; // @[Mux.scala 31:69:@43748.4]
  wire [15:0] _T_100689; // @[Mux.scala 31:69:@43749.4]
  wire [15:0] _T_100690; // @[Mux.scala 31:69:@43750.4]
  wire [15:0] _T_100691; // @[Mux.scala 31:69:@43751.4]
  wire [15:0] _T_100692; // @[Mux.scala 31:69:@43752.4]
  wire [15:0] _T_100693; // @[Mux.scala 31:69:@43753.4]
  wire [15:0] _T_100694; // @[Mux.scala 31:69:@43754.4]
  wire [15:0] _T_100695; // @[Mux.scala 31:69:@43755.4]
  wire [15:0] _T_100696; // @[Mux.scala 31:69:@43756.4]
  wire [15:0] _T_100697; // @[Mux.scala 31:69:@43757.4]
  wire [15:0] _T_100698; // @[Mux.scala 31:69:@43758.4]
  wire [15:0] _T_100699; // @[Mux.scala 31:69:@43759.4]
  wire [15:0] _T_100700; // @[Mux.scala 31:69:@43760.4]
  wire [15:0] _T_100701; // @[Mux.scala 31:69:@43761.4]
  wire [15:0] _T_100702; // @[Mux.scala 31:69:@43762.4]
  wire [15:0] _T_100703; // @[Mux.scala 31:69:@43763.4]
  wire  _T_100704; // @[OneHot.scala 66:30:@43764.4]
  wire  _T_100705; // @[OneHot.scala 66:30:@43765.4]
  wire  _T_100706; // @[OneHot.scala 66:30:@43766.4]
  wire  _T_100707; // @[OneHot.scala 66:30:@43767.4]
  wire  _T_100708; // @[OneHot.scala 66:30:@43768.4]
  wire  _T_100709; // @[OneHot.scala 66:30:@43769.4]
  wire  _T_100710; // @[OneHot.scala 66:30:@43770.4]
  wire  _T_100711; // @[OneHot.scala 66:30:@43771.4]
  wire  _T_100712; // @[OneHot.scala 66:30:@43772.4]
  wire  _T_100713; // @[OneHot.scala 66:30:@43773.4]
  wire  _T_100714; // @[OneHot.scala 66:30:@43774.4]
  wire  _T_100715; // @[OneHot.scala 66:30:@43775.4]
  wire  _T_100716; // @[OneHot.scala 66:30:@43776.4]
  wire  _T_100717; // @[OneHot.scala 66:30:@43777.4]
  wire  _T_100718; // @[OneHot.scala 66:30:@43778.4]
  wire  _T_100719; // @[OneHot.scala 66:30:@43779.4]
  wire [7:0] _T_100784; // @[Mux.scala 19:72:@43803.4]
  wire [15:0] _T_100792; // @[Mux.scala 19:72:@43811.4]
  wire [15:0] _T_100794; // @[Mux.scala 19:72:@43812.4]
  wire [7:0] _T_100801; // @[Mux.scala 19:72:@43819.4]
  wire [15:0] _T_100809; // @[Mux.scala 19:72:@43827.4]
  wire [15:0] _T_100811; // @[Mux.scala 19:72:@43828.4]
  wire [7:0] _T_100818; // @[Mux.scala 19:72:@43835.4]
  wire [15:0] _T_100826; // @[Mux.scala 19:72:@43843.4]
  wire [15:0] _T_100828; // @[Mux.scala 19:72:@43844.4]
  wire [7:0] _T_100835; // @[Mux.scala 19:72:@43851.4]
  wire [15:0] _T_100843; // @[Mux.scala 19:72:@43859.4]
  wire [15:0] _T_100845; // @[Mux.scala 19:72:@43860.4]
  wire [7:0] _T_100852; // @[Mux.scala 19:72:@43867.4]
  wire [15:0] _T_100860; // @[Mux.scala 19:72:@43875.4]
  wire [15:0] _T_100862; // @[Mux.scala 19:72:@43876.4]
  wire [7:0] _T_100869; // @[Mux.scala 19:72:@43883.4]
  wire [15:0] _T_100877; // @[Mux.scala 19:72:@43891.4]
  wire [15:0] _T_100879; // @[Mux.scala 19:72:@43892.4]
  wire [7:0] _T_100886; // @[Mux.scala 19:72:@43899.4]
  wire [15:0] _T_100894; // @[Mux.scala 19:72:@43907.4]
  wire [15:0] _T_100896; // @[Mux.scala 19:72:@43908.4]
  wire [7:0] _T_100903; // @[Mux.scala 19:72:@43915.4]
  wire [15:0] _T_100911; // @[Mux.scala 19:72:@43923.4]
  wire [15:0] _T_100913; // @[Mux.scala 19:72:@43924.4]
  wire [7:0] _T_100920; // @[Mux.scala 19:72:@43931.4]
  wire [15:0] _T_100928; // @[Mux.scala 19:72:@43939.4]
  wire [15:0] _T_100930; // @[Mux.scala 19:72:@43940.4]
  wire [7:0] _T_100937; // @[Mux.scala 19:72:@43947.4]
  wire [15:0] _T_100945; // @[Mux.scala 19:72:@43955.4]
  wire [15:0] _T_100947; // @[Mux.scala 19:72:@43956.4]
  wire [7:0] _T_100954; // @[Mux.scala 19:72:@43963.4]
  wire [15:0] _T_100962; // @[Mux.scala 19:72:@43971.4]
  wire [15:0] _T_100964; // @[Mux.scala 19:72:@43972.4]
  wire [7:0] _T_100971; // @[Mux.scala 19:72:@43979.4]
  wire [15:0] _T_100979; // @[Mux.scala 19:72:@43987.4]
  wire [15:0] _T_100981; // @[Mux.scala 19:72:@43988.4]
  wire [7:0] _T_100988; // @[Mux.scala 19:72:@43995.4]
  wire [15:0] _T_100996; // @[Mux.scala 19:72:@44003.4]
  wire [15:0] _T_100998; // @[Mux.scala 19:72:@44004.4]
  wire [7:0] _T_101005; // @[Mux.scala 19:72:@44011.4]
  wire [15:0] _T_101013; // @[Mux.scala 19:72:@44019.4]
  wire [15:0] _T_101015; // @[Mux.scala 19:72:@44020.4]
  wire [7:0] _T_101022; // @[Mux.scala 19:72:@44027.4]
  wire [15:0] _T_101030; // @[Mux.scala 19:72:@44035.4]
  wire [15:0] _T_101032; // @[Mux.scala 19:72:@44036.4]
  wire [7:0] _T_101039; // @[Mux.scala 19:72:@44043.4]
  wire [15:0] _T_101047; // @[Mux.scala 19:72:@44051.4]
  wire [15:0] _T_101049; // @[Mux.scala 19:72:@44052.4]
  wire [15:0] _T_101050; // @[Mux.scala 19:72:@44053.4]
  wire [15:0] _T_101051; // @[Mux.scala 19:72:@44054.4]
  wire [15:0] _T_101052; // @[Mux.scala 19:72:@44055.4]
  wire [15:0] _T_101053; // @[Mux.scala 19:72:@44056.4]
  wire [15:0] _T_101054; // @[Mux.scala 19:72:@44057.4]
  wire [15:0] _T_101055; // @[Mux.scala 19:72:@44058.4]
  wire [15:0] _T_101056; // @[Mux.scala 19:72:@44059.4]
  wire [15:0] _T_101057; // @[Mux.scala 19:72:@44060.4]
  wire [15:0] _T_101058; // @[Mux.scala 19:72:@44061.4]
  wire [15:0] _T_101059; // @[Mux.scala 19:72:@44062.4]
  wire [15:0] _T_101060; // @[Mux.scala 19:72:@44063.4]
  wire [15:0] _T_101061; // @[Mux.scala 19:72:@44064.4]
  wire [15:0] _T_101062; // @[Mux.scala 19:72:@44065.4]
  wire [15:0] _T_101063; // @[Mux.scala 19:72:@44066.4]
  wire [15:0] _T_101064; // @[Mux.scala 19:72:@44067.4]
  wire  outputPriorityPorts_1_0; // @[Mux.scala 19:72:@44071.4]
  wire  outputPriorityPorts_1_1; // @[Mux.scala 19:72:@44073.4]
  wire  outputPriorityPorts_1_2; // @[Mux.scala 19:72:@44075.4]
  wire  outputPriorityPorts_1_3; // @[Mux.scala 19:72:@44077.4]
  wire  outputPriorityPorts_1_4; // @[Mux.scala 19:72:@44079.4]
  wire  outputPriorityPorts_1_5; // @[Mux.scala 19:72:@44081.4]
  wire  outputPriorityPorts_1_6; // @[Mux.scala 19:72:@44083.4]
  wire  outputPriorityPorts_1_7; // @[Mux.scala 19:72:@44085.4]
  wire  outputPriorityPorts_1_8; // @[Mux.scala 19:72:@44087.4]
  wire  outputPriorityPorts_1_9; // @[Mux.scala 19:72:@44089.4]
  wire  outputPriorityPorts_1_10; // @[Mux.scala 19:72:@44091.4]
  wire  outputPriorityPorts_1_11; // @[Mux.scala 19:72:@44093.4]
  wire  outputPriorityPorts_1_12; // @[Mux.scala 19:72:@44095.4]
  wire  outputPriorityPorts_1_13; // @[Mux.scala 19:72:@44097.4]
  wire  outputPriorityPorts_1_14; // @[Mux.scala 19:72:@44099.4]
  wire  outputPriorityPorts_1_15; // @[Mux.scala 19:72:@44101.4]
  wire  _T_101207; // @[LoadQueue.scala 313:47:@44123.6]
  wire  _T_101208; // @[LoadQueue.scala 313:47:@44124.6]
  wire  _T_101219; // @[LoadQueue.scala 314:26:@44129.6]
  wire [1:0] _T_101220; // @[OneHot.scala 18:45:@44131.8]
  wire  _T_101221; // @[CircuitMath.scala 30:8:@44132.8]
  wire [31:0] _GEN_2115; // @[LoadQueue.scala 315:29:@44133.8]
  wire [31:0] _GEN_2116; // @[LoadQueue.scala 314:36:@44130.6]
  wire  _GEN_2117; // @[LoadQueue.scala 314:36:@44130.6]
  wire  _GEN_2118; // @[LoadQueue.scala 308:34:@44119.4]
  wire [31:0] _GEN_2119; // @[LoadQueue.scala 308:34:@44119.4]
  wire  _T_101225; // @[LoadQueue.scala 313:47:@44141.6]
  wire  _T_101226; // @[LoadQueue.scala 313:47:@44142.6]
  wire  _T_101237; // @[LoadQueue.scala 314:26:@44147.6]
  wire [1:0] _T_101238; // @[OneHot.scala 18:45:@44149.8]
  wire  _T_101239; // @[CircuitMath.scala 30:8:@44150.8]
  wire [31:0] _GEN_2121; // @[LoadQueue.scala 315:29:@44151.8]
  wire [31:0] _GEN_2122; // @[LoadQueue.scala 314:36:@44148.6]
  wire  _GEN_2123; // @[LoadQueue.scala 314:36:@44148.6]
  wire  _GEN_2124; // @[LoadQueue.scala 308:34:@44137.4]
  wire [31:0] _GEN_2125; // @[LoadQueue.scala 308:34:@44137.4]
  wire  _T_101243; // @[LoadQueue.scala 313:47:@44159.6]
  wire  _T_101244; // @[LoadQueue.scala 313:47:@44160.6]
  wire  _T_101255; // @[LoadQueue.scala 314:26:@44165.6]
  wire [1:0] _T_101256; // @[OneHot.scala 18:45:@44167.8]
  wire  _T_101257; // @[CircuitMath.scala 30:8:@44168.8]
  wire [31:0] _GEN_2127; // @[LoadQueue.scala 315:29:@44169.8]
  wire [31:0] _GEN_2128; // @[LoadQueue.scala 314:36:@44166.6]
  wire  _GEN_2129; // @[LoadQueue.scala 314:36:@44166.6]
  wire  _GEN_2130; // @[LoadQueue.scala 308:34:@44155.4]
  wire [31:0] _GEN_2131; // @[LoadQueue.scala 308:34:@44155.4]
  wire  _T_101261; // @[LoadQueue.scala 313:47:@44177.6]
  wire  _T_101262; // @[LoadQueue.scala 313:47:@44178.6]
  wire  _T_101273; // @[LoadQueue.scala 314:26:@44183.6]
  wire [1:0] _T_101274; // @[OneHot.scala 18:45:@44185.8]
  wire  _T_101275; // @[CircuitMath.scala 30:8:@44186.8]
  wire [31:0] _GEN_2133; // @[LoadQueue.scala 315:29:@44187.8]
  wire [31:0] _GEN_2134; // @[LoadQueue.scala 314:36:@44184.6]
  wire  _GEN_2135; // @[LoadQueue.scala 314:36:@44184.6]
  wire  _GEN_2136; // @[LoadQueue.scala 308:34:@44173.4]
  wire [31:0] _GEN_2137; // @[LoadQueue.scala 308:34:@44173.4]
  wire  _T_101279; // @[LoadQueue.scala 313:47:@44195.6]
  wire  _T_101280; // @[LoadQueue.scala 313:47:@44196.6]
  wire  _T_101291; // @[LoadQueue.scala 314:26:@44201.6]
  wire [1:0] _T_101292; // @[OneHot.scala 18:45:@44203.8]
  wire  _T_101293; // @[CircuitMath.scala 30:8:@44204.8]
  wire [31:0] _GEN_2139; // @[LoadQueue.scala 315:29:@44205.8]
  wire [31:0] _GEN_2140; // @[LoadQueue.scala 314:36:@44202.6]
  wire  _GEN_2141; // @[LoadQueue.scala 314:36:@44202.6]
  wire  _GEN_2142; // @[LoadQueue.scala 308:34:@44191.4]
  wire [31:0] _GEN_2143; // @[LoadQueue.scala 308:34:@44191.4]
  wire  _T_101297; // @[LoadQueue.scala 313:47:@44213.6]
  wire  _T_101298; // @[LoadQueue.scala 313:47:@44214.6]
  wire  _T_101309; // @[LoadQueue.scala 314:26:@44219.6]
  wire [1:0] _T_101310; // @[OneHot.scala 18:45:@44221.8]
  wire  _T_101311; // @[CircuitMath.scala 30:8:@44222.8]
  wire [31:0] _GEN_2145; // @[LoadQueue.scala 315:29:@44223.8]
  wire [31:0] _GEN_2146; // @[LoadQueue.scala 314:36:@44220.6]
  wire  _GEN_2147; // @[LoadQueue.scala 314:36:@44220.6]
  wire  _GEN_2148; // @[LoadQueue.scala 308:34:@44209.4]
  wire [31:0] _GEN_2149; // @[LoadQueue.scala 308:34:@44209.4]
  wire  _T_101315; // @[LoadQueue.scala 313:47:@44231.6]
  wire  _T_101316; // @[LoadQueue.scala 313:47:@44232.6]
  wire  _T_101327; // @[LoadQueue.scala 314:26:@44237.6]
  wire [1:0] _T_101328; // @[OneHot.scala 18:45:@44239.8]
  wire  _T_101329; // @[CircuitMath.scala 30:8:@44240.8]
  wire [31:0] _GEN_2151; // @[LoadQueue.scala 315:29:@44241.8]
  wire [31:0] _GEN_2152; // @[LoadQueue.scala 314:36:@44238.6]
  wire  _GEN_2153; // @[LoadQueue.scala 314:36:@44238.6]
  wire  _GEN_2154; // @[LoadQueue.scala 308:34:@44227.4]
  wire [31:0] _GEN_2155; // @[LoadQueue.scala 308:34:@44227.4]
  wire  _T_101333; // @[LoadQueue.scala 313:47:@44249.6]
  wire  _T_101334; // @[LoadQueue.scala 313:47:@44250.6]
  wire  _T_101345; // @[LoadQueue.scala 314:26:@44255.6]
  wire [1:0] _T_101346; // @[OneHot.scala 18:45:@44257.8]
  wire  _T_101347; // @[CircuitMath.scala 30:8:@44258.8]
  wire [31:0] _GEN_2157; // @[LoadQueue.scala 315:29:@44259.8]
  wire [31:0] _GEN_2158; // @[LoadQueue.scala 314:36:@44256.6]
  wire  _GEN_2159; // @[LoadQueue.scala 314:36:@44256.6]
  wire  _GEN_2160; // @[LoadQueue.scala 308:34:@44245.4]
  wire [31:0] _GEN_2161; // @[LoadQueue.scala 308:34:@44245.4]
  wire  _T_101351; // @[LoadQueue.scala 313:47:@44267.6]
  wire  _T_101352; // @[LoadQueue.scala 313:47:@44268.6]
  wire  _T_101363; // @[LoadQueue.scala 314:26:@44273.6]
  wire [1:0] _T_101364; // @[OneHot.scala 18:45:@44275.8]
  wire  _T_101365; // @[CircuitMath.scala 30:8:@44276.8]
  wire [31:0] _GEN_2163; // @[LoadQueue.scala 315:29:@44277.8]
  wire [31:0] _GEN_2164; // @[LoadQueue.scala 314:36:@44274.6]
  wire  _GEN_2165; // @[LoadQueue.scala 314:36:@44274.6]
  wire  _GEN_2166; // @[LoadQueue.scala 308:34:@44263.4]
  wire [31:0] _GEN_2167; // @[LoadQueue.scala 308:34:@44263.4]
  wire  _T_101369; // @[LoadQueue.scala 313:47:@44285.6]
  wire  _T_101370; // @[LoadQueue.scala 313:47:@44286.6]
  wire  _T_101381; // @[LoadQueue.scala 314:26:@44291.6]
  wire [1:0] _T_101382; // @[OneHot.scala 18:45:@44293.8]
  wire  _T_101383; // @[CircuitMath.scala 30:8:@44294.8]
  wire [31:0] _GEN_2169; // @[LoadQueue.scala 315:29:@44295.8]
  wire [31:0] _GEN_2170; // @[LoadQueue.scala 314:36:@44292.6]
  wire  _GEN_2171; // @[LoadQueue.scala 314:36:@44292.6]
  wire  _GEN_2172; // @[LoadQueue.scala 308:34:@44281.4]
  wire [31:0] _GEN_2173; // @[LoadQueue.scala 308:34:@44281.4]
  wire  _T_101387; // @[LoadQueue.scala 313:47:@44303.6]
  wire  _T_101388; // @[LoadQueue.scala 313:47:@44304.6]
  wire  _T_101399; // @[LoadQueue.scala 314:26:@44309.6]
  wire [1:0] _T_101400; // @[OneHot.scala 18:45:@44311.8]
  wire  _T_101401; // @[CircuitMath.scala 30:8:@44312.8]
  wire [31:0] _GEN_2175; // @[LoadQueue.scala 315:29:@44313.8]
  wire [31:0] _GEN_2176; // @[LoadQueue.scala 314:36:@44310.6]
  wire  _GEN_2177; // @[LoadQueue.scala 314:36:@44310.6]
  wire  _GEN_2178; // @[LoadQueue.scala 308:34:@44299.4]
  wire [31:0] _GEN_2179; // @[LoadQueue.scala 308:34:@44299.4]
  wire  _T_101405; // @[LoadQueue.scala 313:47:@44321.6]
  wire  _T_101406; // @[LoadQueue.scala 313:47:@44322.6]
  wire  _T_101417; // @[LoadQueue.scala 314:26:@44327.6]
  wire [1:0] _T_101418; // @[OneHot.scala 18:45:@44329.8]
  wire  _T_101419; // @[CircuitMath.scala 30:8:@44330.8]
  wire [31:0] _GEN_2181; // @[LoadQueue.scala 315:29:@44331.8]
  wire [31:0] _GEN_2182; // @[LoadQueue.scala 314:36:@44328.6]
  wire  _GEN_2183; // @[LoadQueue.scala 314:36:@44328.6]
  wire  _GEN_2184; // @[LoadQueue.scala 308:34:@44317.4]
  wire [31:0] _GEN_2185; // @[LoadQueue.scala 308:34:@44317.4]
  wire  _T_101423; // @[LoadQueue.scala 313:47:@44339.6]
  wire  _T_101424; // @[LoadQueue.scala 313:47:@44340.6]
  wire  _T_101435; // @[LoadQueue.scala 314:26:@44345.6]
  wire [1:0] _T_101436; // @[OneHot.scala 18:45:@44347.8]
  wire  _T_101437; // @[CircuitMath.scala 30:8:@44348.8]
  wire [31:0] _GEN_2187; // @[LoadQueue.scala 315:29:@44349.8]
  wire [31:0] _GEN_2188; // @[LoadQueue.scala 314:36:@44346.6]
  wire  _GEN_2189; // @[LoadQueue.scala 314:36:@44346.6]
  wire  _GEN_2190; // @[LoadQueue.scala 308:34:@44335.4]
  wire [31:0] _GEN_2191; // @[LoadQueue.scala 308:34:@44335.4]
  wire  _T_101441; // @[LoadQueue.scala 313:47:@44357.6]
  wire  _T_101442; // @[LoadQueue.scala 313:47:@44358.6]
  wire  _T_101453; // @[LoadQueue.scala 314:26:@44363.6]
  wire [1:0] _T_101454; // @[OneHot.scala 18:45:@44365.8]
  wire  _T_101455; // @[CircuitMath.scala 30:8:@44366.8]
  wire [31:0] _GEN_2193; // @[LoadQueue.scala 315:29:@44367.8]
  wire [31:0] _GEN_2194; // @[LoadQueue.scala 314:36:@44364.6]
  wire  _GEN_2195; // @[LoadQueue.scala 314:36:@44364.6]
  wire  _GEN_2196; // @[LoadQueue.scala 308:34:@44353.4]
  wire [31:0] _GEN_2197; // @[LoadQueue.scala 308:34:@44353.4]
  wire  _T_101459; // @[LoadQueue.scala 313:47:@44375.6]
  wire  _T_101460; // @[LoadQueue.scala 313:47:@44376.6]
  wire  _T_101471; // @[LoadQueue.scala 314:26:@44381.6]
  wire [1:0] _T_101472; // @[OneHot.scala 18:45:@44383.8]
  wire  _T_101473; // @[CircuitMath.scala 30:8:@44384.8]
  wire [31:0] _GEN_2199; // @[LoadQueue.scala 315:29:@44385.8]
  wire [31:0] _GEN_2200; // @[LoadQueue.scala 314:36:@44382.6]
  wire  _GEN_2201; // @[LoadQueue.scala 314:36:@44382.6]
  wire  _GEN_2202; // @[LoadQueue.scala 308:34:@44371.4]
  wire [31:0] _GEN_2203; // @[LoadQueue.scala 308:34:@44371.4]
  wire  _T_101477; // @[LoadQueue.scala 313:47:@44393.6]
  wire  _T_101478; // @[LoadQueue.scala 313:47:@44394.6]
  wire  _T_101489; // @[LoadQueue.scala 314:26:@44399.6]
  wire [1:0] _T_101490; // @[OneHot.scala 18:45:@44401.8]
  wire  _T_101491; // @[CircuitMath.scala 30:8:@44402.8]
  wire [31:0] _GEN_2205; // @[LoadQueue.scala 315:29:@44403.8]
  wire [31:0] _GEN_2206; // @[LoadQueue.scala 314:36:@44400.6]
  wire  _GEN_2207; // @[LoadQueue.scala 314:36:@44400.6]
  wire  _GEN_2208; // @[LoadQueue.scala 308:34:@44389.4]
  wire [31:0] _GEN_2209; // @[LoadQueue.scala 308:34:@44389.4]
  wire  _T_101515; // @[LoadQueue.scala 326:108:@44408.4]
  wire  _T_101517; // @[LoadQueue.scala 327:34:@44409.4]
  wire  _T_101518; // @[LoadQueue.scala 327:31:@44410.4]
  wire  _T_101519; // @[LoadQueue.scala 327:63:@44411.4]
  wire  _T_101520; // @[LoadQueue.scala 326:108:@44412.4]
  wire  _T_101523; // @[LoadQueue.scala 327:31:@44414.4]
  wire  _T_101524; // @[LoadQueue.scala 327:63:@44415.4]
  wire  loadCompleting_0; // @[LoadQueue.scala 328:51:@44420.4]
  wire  _T_101536; // @[LoadQueue.scala 326:108:@44422.4]
  wire  _T_101538; // @[LoadQueue.scala 327:34:@44423.4]
  wire  _T_101539; // @[LoadQueue.scala 327:31:@44424.4]
  wire  _T_101540; // @[LoadQueue.scala 327:63:@44425.4]
  wire  _T_101541; // @[LoadQueue.scala 326:108:@44426.4]
  wire  _T_101544; // @[LoadQueue.scala 327:31:@44428.4]
  wire  _T_101545; // @[LoadQueue.scala 327:63:@44429.4]
  wire  loadCompleting_1; // @[LoadQueue.scala 328:51:@44434.4]
  wire  _T_101557; // @[LoadQueue.scala 326:108:@44436.4]
  wire  _T_101559; // @[LoadQueue.scala 327:34:@44437.4]
  wire  _T_101560; // @[LoadQueue.scala 327:31:@44438.4]
  wire  _T_101561; // @[LoadQueue.scala 327:63:@44439.4]
  wire  _T_101562; // @[LoadQueue.scala 326:108:@44440.4]
  wire  _T_101565; // @[LoadQueue.scala 327:31:@44442.4]
  wire  _T_101566; // @[LoadQueue.scala 327:63:@44443.4]
  wire  loadCompleting_2; // @[LoadQueue.scala 328:51:@44448.4]
  wire  _T_101578; // @[LoadQueue.scala 326:108:@44450.4]
  wire  _T_101580; // @[LoadQueue.scala 327:34:@44451.4]
  wire  _T_101581; // @[LoadQueue.scala 327:31:@44452.4]
  wire  _T_101582; // @[LoadQueue.scala 327:63:@44453.4]
  wire  _T_101583; // @[LoadQueue.scala 326:108:@44454.4]
  wire  _T_101586; // @[LoadQueue.scala 327:31:@44456.4]
  wire  _T_101587; // @[LoadQueue.scala 327:63:@44457.4]
  wire  loadCompleting_3; // @[LoadQueue.scala 328:51:@44462.4]
  wire  _T_101599; // @[LoadQueue.scala 326:108:@44464.4]
  wire  _T_101601; // @[LoadQueue.scala 327:34:@44465.4]
  wire  _T_101602; // @[LoadQueue.scala 327:31:@44466.4]
  wire  _T_101603; // @[LoadQueue.scala 327:63:@44467.4]
  wire  _T_101604; // @[LoadQueue.scala 326:108:@44468.4]
  wire  _T_101607; // @[LoadQueue.scala 327:31:@44470.4]
  wire  _T_101608; // @[LoadQueue.scala 327:63:@44471.4]
  wire  loadCompleting_4; // @[LoadQueue.scala 328:51:@44476.4]
  wire  _T_101620; // @[LoadQueue.scala 326:108:@44478.4]
  wire  _T_101622; // @[LoadQueue.scala 327:34:@44479.4]
  wire  _T_101623; // @[LoadQueue.scala 327:31:@44480.4]
  wire  _T_101624; // @[LoadQueue.scala 327:63:@44481.4]
  wire  _T_101625; // @[LoadQueue.scala 326:108:@44482.4]
  wire  _T_101628; // @[LoadQueue.scala 327:31:@44484.4]
  wire  _T_101629; // @[LoadQueue.scala 327:63:@44485.4]
  wire  loadCompleting_5; // @[LoadQueue.scala 328:51:@44490.4]
  wire  _T_101641; // @[LoadQueue.scala 326:108:@44492.4]
  wire  _T_101643; // @[LoadQueue.scala 327:34:@44493.4]
  wire  _T_101644; // @[LoadQueue.scala 327:31:@44494.4]
  wire  _T_101645; // @[LoadQueue.scala 327:63:@44495.4]
  wire  _T_101646; // @[LoadQueue.scala 326:108:@44496.4]
  wire  _T_101649; // @[LoadQueue.scala 327:31:@44498.4]
  wire  _T_101650; // @[LoadQueue.scala 327:63:@44499.4]
  wire  loadCompleting_6; // @[LoadQueue.scala 328:51:@44504.4]
  wire  _T_101662; // @[LoadQueue.scala 326:108:@44506.4]
  wire  _T_101664; // @[LoadQueue.scala 327:34:@44507.4]
  wire  _T_101665; // @[LoadQueue.scala 327:31:@44508.4]
  wire  _T_101666; // @[LoadQueue.scala 327:63:@44509.4]
  wire  _T_101667; // @[LoadQueue.scala 326:108:@44510.4]
  wire  _T_101670; // @[LoadQueue.scala 327:31:@44512.4]
  wire  _T_101671; // @[LoadQueue.scala 327:63:@44513.4]
  wire  loadCompleting_7; // @[LoadQueue.scala 328:51:@44518.4]
  wire  _T_101683; // @[LoadQueue.scala 326:108:@44520.4]
  wire  _T_101685; // @[LoadQueue.scala 327:34:@44521.4]
  wire  _T_101686; // @[LoadQueue.scala 327:31:@44522.4]
  wire  _T_101687; // @[LoadQueue.scala 327:63:@44523.4]
  wire  _T_101688; // @[LoadQueue.scala 326:108:@44524.4]
  wire  _T_101691; // @[LoadQueue.scala 327:31:@44526.4]
  wire  _T_101692; // @[LoadQueue.scala 327:63:@44527.4]
  wire  loadCompleting_8; // @[LoadQueue.scala 328:51:@44532.4]
  wire  _T_101704; // @[LoadQueue.scala 326:108:@44534.4]
  wire  _T_101706; // @[LoadQueue.scala 327:34:@44535.4]
  wire  _T_101707; // @[LoadQueue.scala 327:31:@44536.4]
  wire  _T_101708; // @[LoadQueue.scala 327:63:@44537.4]
  wire  _T_101709; // @[LoadQueue.scala 326:108:@44538.4]
  wire  _T_101712; // @[LoadQueue.scala 327:31:@44540.4]
  wire  _T_101713; // @[LoadQueue.scala 327:63:@44541.4]
  wire  loadCompleting_9; // @[LoadQueue.scala 328:51:@44546.4]
  wire  _T_101725; // @[LoadQueue.scala 326:108:@44548.4]
  wire  _T_101727; // @[LoadQueue.scala 327:34:@44549.4]
  wire  _T_101728; // @[LoadQueue.scala 327:31:@44550.4]
  wire  _T_101729; // @[LoadQueue.scala 327:63:@44551.4]
  wire  _T_101730; // @[LoadQueue.scala 326:108:@44552.4]
  wire  _T_101733; // @[LoadQueue.scala 327:31:@44554.4]
  wire  _T_101734; // @[LoadQueue.scala 327:63:@44555.4]
  wire  loadCompleting_10; // @[LoadQueue.scala 328:51:@44560.4]
  wire  _T_101746; // @[LoadQueue.scala 326:108:@44562.4]
  wire  _T_101748; // @[LoadQueue.scala 327:34:@44563.4]
  wire  _T_101749; // @[LoadQueue.scala 327:31:@44564.4]
  wire  _T_101750; // @[LoadQueue.scala 327:63:@44565.4]
  wire  _T_101751; // @[LoadQueue.scala 326:108:@44566.4]
  wire  _T_101754; // @[LoadQueue.scala 327:31:@44568.4]
  wire  _T_101755; // @[LoadQueue.scala 327:63:@44569.4]
  wire  loadCompleting_11; // @[LoadQueue.scala 328:51:@44574.4]
  wire  _T_101767; // @[LoadQueue.scala 326:108:@44576.4]
  wire  _T_101769; // @[LoadQueue.scala 327:34:@44577.4]
  wire  _T_101770; // @[LoadQueue.scala 327:31:@44578.4]
  wire  _T_101771; // @[LoadQueue.scala 327:63:@44579.4]
  wire  _T_101772; // @[LoadQueue.scala 326:108:@44580.4]
  wire  _T_101775; // @[LoadQueue.scala 327:31:@44582.4]
  wire  _T_101776; // @[LoadQueue.scala 327:63:@44583.4]
  wire  loadCompleting_12; // @[LoadQueue.scala 328:51:@44588.4]
  wire  _T_101788; // @[LoadQueue.scala 326:108:@44590.4]
  wire  _T_101790; // @[LoadQueue.scala 327:34:@44591.4]
  wire  _T_101791; // @[LoadQueue.scala 327:31:@44592.4]
  wire  _T_101792; // @[LoadQueue.scala 327:63:@44593.4]
  wire  _T_101793; // @[LoadQueue.scala 326:108:@44594.4]
  wire  _T_101796; // @[LoadQueue.scala 327:31:@44596.4]
  wire  _T_101797; // @[LoadQueue.scala 327:63:@44597.4]
  wire  loadCompleting_13; // @[LoadQueue.scala 328:51:@44602.4]
  wire  _T_101809; // @[LoadQueue.scala 326:108:@44604.4]
  wire  _T_101811; // @[LoadQueue.scala 327:34:@44605.4]
  wire  _T_101812; // @[LoadQueue.scala 327:31:@44606.4]
  wire  _T_101813; // @[LoadQueue.scala 327:63:@44607.4]
  wire  _T_101814; // @[LoadQueue.scala 326:108:@44608.4]
  wire  _T_101817; // @[LoadQueue.scala 327:31:@44610.4]
  wire  _T_101818; // @[LoadQueue.scala 327:63:@44611.4]
  wire  loadCompleting_14; // @[LoadQueue.scala 328:51:@44616.4]
  wire  _T_101830; // @[LoadQueue.scala 326:108:@44618.4]
  wire  _T_101832; // @[LoadQueue.scala 327:34:@44619.4]
  wire  _T_101833; // @[LoadQueue.scala 327:31:@44620.4]
  wire  _T_101834; // @[LoadQueue.scala 327:63:@44621.4]
  wire  _T_101835; // @[LoadQueue.scala 326:108:@44622.4]
  wire  _T_101838; // @[LoadQueue.scala 327:31:@44624.4]
  wire  _T_101839; // @[LoadQueue.scala 327:63:@44625.4]
  wire  loadCompleting_15; // @[LoadQueue.scala 328:51:@44630.4]
  wire  _GEN_2210; // @[LoadQueue.scala 337:46:@44636.6]
  wire  _GEN_2211; // @[LoadQueue.scala 335:34:@44632.4]
  wire  _GEN_2212; // @[LoadQueue.scala 337:46:@44643.6]
  wire  _GEN_2213; // @[LoadQueue.scala 335:34:@44639.4]
  wire  _GEN_2214; // @[LoadQueue.scala 337:46:@44650.6]
  wire  _GEN_2215; // @[LoadQueue.scala 335:34:@44646.4]
  wire  _GEN_2216; // @[LoadQueue.scala 337:46:@44657.6]
  wire  _GEN_2217; // @[LoadQueue.scala 335:34:@44653.4]
  wire  _GEN_2218; // @[LoadQueue.scala 337:46:@44664.6]
  wire  _GEN_2219; // @[LoadQueue.scala 335:34:@44660.4]
  wire  _GEN_2220; // @[LoadQueue.scala 337:46:@44671.6]
  wire  _GEN_2221; // @[LoadQueue.scala 335:34:@44667.4]
  wire  _GEN_2222; // @[LoadQueue.scala 337:46:@44678.6]
  wire  _GEN_2223; // @[LoadQueue.scala 335:34:@44674.4]
  wire  _GEN_2224; // @[LoadQueue.scala 337:46:@44685.6]
  wire  _GEN_2225; // @[LoadQueue.scala 335:34:@44681.4]
  wire  _GEN_2226; // @[LoadQueue.scala 337:46:@44692.6]
  wire  _GEN_2227; // @[LoadQueue.scala 335:34:@44688.4]
  wire  _GEN_2228; // @[LoadQueue.scala 337:46:@44699.6]
  wire  _GEN_2229; // @[LoadQueue.scala 335:34:@44695.4]
  wire  _GEN_2230; // @[LoadQueue.scala 337:46:@44706.6]
  wire  _GEN_2231; // @[LoadQueue.scala 335:34:@44702.4]
  wire  _GEN_2232; // @[LoadQueue.scala 337:46:@44713.6]
  wire  _GEN_2233; // @[LoadQueue.scala 335:34:@44709.4]
  wire  _GEN_2234; // @[LoadQueue.scala 337:46:@44720.6]
  wire  _GEN_2235; // @[LoadQueue.scala 335:34:@44716.4]
  wire  _GEN_2236; // @[LoadQueue.scala 337:46:@44727.6]
  wire  _GEN_2237; // @[LoadQueue.scala 335:34:@44723.4]
  wire  _GEN_2238; // @[LoadQueue.scala 337:46:@44734.6]
  wire  _GEN_2239; // @[LoadQueue.scala 335:34:@44730.4]
  wire  _GEN_2240; // @[LoadQueue.scala 337:46:@44741.6]
  wire  _GEN_2241; // @[LoadQueue.scala 335:34:@44737.4]
  wire  _T_101971; // @[LoadQueue.scala 348:24:@44810.4]
  wire  _T_101972; // @[LoadQueue.scala 348:24:@44811.4]
  wire  _T_101973; // @[LoadQueue.scala 348:24:@44812.4]
  wire  _T_101974; // @[LoadQueue.scala 348:24:@44813.4]
  wire  _T_101975; // @[LoadQueue.scala 348:24:@44814.4]
  wire  _T_101976; // @[LoadQueue.scala 348:24:@44815.4]
  wire  _T_101977; // @[LoadQueue.scala 348:24:@44816.4]
  wire  _T_101978; // @[LoadQueue.scala 348:24:@44817.4]
  wire  _T_101979; // @[LoadQueue.scala 348:24:@44818.4]
  wire  _T_101980; // @[LoadQueue.scala 348:24:@44819.4]
  wire  _T_101981; // @[LoadQueue.scala 348:24:@44820.4]
  wire  _T_101982; // @[LoadQueue.scala 348:24:@44821.4]
  wire  _T_101983; // @[LoadQueue.scala 348:24:@44822.4]
  wire  _T_101984; // @[LoadQueue.scala 348:24:@44823.4]
  wire  _T_101985; // @[LoadQueue.scala 348:24:@44824.4]
  wire [3:0] _T_102002; // @[Mux.scala 31:69:@44826.6]
  wire [3:0] _T_102003; // @[Mux.scala 31:69:@44827.6]
  wire [3:0] _T_102004; // @[Mux.scala 31:69:@44828.6]
  wire [3:0] _T_102005; // @[Mux.scala 31:69:@44829.6]
  wire [3:0] _T_102006; // @[Mux.scala 31:69:@44830.6]
  wire [3:0] _T_102007; // @[Mux.scala 31:69:@44831.6]
  wire [3:0] _T_102008; // @[Mux.scala 31:69:@44832.6]
  wire [3:0] _T_102009; // @[Mux.scala 31:69:@44833.6]
  wire [3:0] _T_102010; // @[Mux.scala 31:69:@44834.6]
  wire [3:0] _T_102011; // @[Mux.scala 31:69:@44835.6]
  wire [3:0] _T_102012; // @[Mux.scala 31:69:@44836.6]
  wire [3:0] _T_102013; // @[Mux.scala 31:69:@44837.6]
  wire [3:0] _T_102014; // @[Mux.scala 31:69:@44838.6]
  wire [3:0] _T_102015; // @[Mux.scala 31:69:@44839.6]
  wire [3:0] _T_102016; // @[Mux.scala 31:69:@44840.6]
  wire [31:0] _GEN_2243; // @[LoadQueue.scala 349:37:@44841.6]
  wire [31:0] _GEN_2244; // @[LoadQueue.scala 349:37:@44841.6]
  wire [31:0] _GEN_2245; // @[LoadQueue.scala 349:37:@44841.6]
  wire [31:0] _GEN_2246; // @[LoadQueue.scala 349:37:@44841.6]
  wire [31:0] _GEN_2247; // @[LoadQueue.scala 349:37:@44841.6]
  wire [31:0] _GEN_2248; // @[LoadQueue.scala 349:37:@44841.6]
  wire [31:0] _GEN_2249; // @[LoadQueue.scala 349:37:@44841.6]
  wire [31:0] _GEN_2250; // @[LoadQueue.scala 349:37:@44841.6]
  wire [31:0] _GEN_2251; // @[LoadQueue.scala 349:37:@44841.6]
  wire [31:0] _GEN_2252; // @[LoadQueue.scala 349:37:@44841.6]
  wire [31:0] _GEN_2253; // @[LoadQueue.scala 349:37:@44841.6]
  wire [31:0] _GEN_2254; // @[LoadQueue.scala 349:37:@44841.6]
  wire [31:0] _GEN_2255; // @[LoadQueue.scala 349:37:@44841.6]
  wire [31:0] _GEN_2256; // @[LoadQueue.scala 349:37:@44841.6]
  wire [31:0] _GEN_2257; // @[LoadQueue.scala 349:37:@44841.6]
  wire  _T_102111; // @[LoadQueue.scala 348:24:@44914.4]
  wire  _T_102112; // @[LoadQueue.scala 348:24:@44915.4]
  wire  _T_102113; // @[LoadQueue.scala 348:24:@44916.4]
  wire  _T_102114; // @[LoadQueue.scala 348:24:@44917.4]
  wire  _T_102115; // @[LoadQueue.scala 348:24:@44918.4]
  wire  _T_102116; // @[LoadQueue.scala 348:24:@44919.4]
  wire  _T_102117; // @[LoadQueue.scala 348:24:@44920.4]
  wire  _T_102118; // @[LoadQueue.scala 348:24:@44921.4]
  wire  _T_102119; // @[LoadQueue.scala 348:24:@44922.4]
  wire  _T_102120; // @[LoadQueue.scala 348:24:@44923.4]
  wire  _T_102121; // @[LoadQueue.scala 348:24:@44924.4]
  wire  _T_102122; // @[LoadQueue.scala 348:24:@44925.4]
  wire  _T_102123; // @[LoadQueue.scala 348:24:@44926.4]
  wire  _T_102124; // @[LoadQueue.scala 348:24:@44927.4]
  wire  _T_102125; // @[LoadQueue.scala 348:24:@44928.4]
  wire [3:0] _T_102142; // @[Mux.scala 31:69:@44930.6]
  wire [3:0] _T_102143; // @[Mux.scala 31:69:@44931.6]
  wire [3:0] _T_102144; // @[Mux.scala 31:69:@44932.6]
  wire [3:0] _T_102145; // @[Mux.scala 31:69:@44933.6]
  wire [3:0] _T_102146; // @[Mux.scala 31:69:@44934.6]
  wire [3:0] _T_102147; // @[Mux.scala 31:69:@44935.6]
  wire [3:0] _T_102148; // @[Mux.scala 31:69:@44936.6]
  wire [3:0] _T_102149; // @[Mux.scala 31:69:@44937.6]
  wire [3:0] _T_102150; // @[Mux.scala 31:69:@44938.6]
  wire [3:0] _T_102151; // @[Mux.scala 31:69:@44939.6]
  wire [3:0] _T_102152; // @[Mux.scala 31:69:@44940.6]
  wire [3:0] _T_102153; // @[Mux.scala 31:69:@44941.6]
  wire [3:0] _T_102154; // @[Mux.scala 31:69:@44942.6]
  wire [3:0] _T_102155; // @[Mux.scala 31:69:@44943.6]
  wire [3:0] _T_102156; // @[Mux.scala 31:69:@44944.6]
  wire [31:0] _GEN_2261; // @[LoadQueue.scala 349:37:@44945.6]
  wire [31:0] _GEN_2262; // @[LoadQueue.scala 349:37:@44945.6]
  wire [31:0] _GEN_2263; // @[LoadQueue.scala 349:37:@44945.6]
  wire [31:0] _GEN_2264; // @[LoadQueue.scala 349:37:@44945.6]
  wire [31:0] _GEN_2265; // @[LoadQueue.scala 349:37:@44945.6]
  wire [31:0] _GEN_2266; // @[LoadQueue.scala 349:37:@44945.6]
  wire [31:0] _GEN_2267; // @[LoadQueue.scala 349:37:@44945.6]
  wire [31:0] _GEN_2268; // @[LoadQueue.scala 349:37:@44945.6]
  wire [31:0] _GEN_2269; // @[LoadQueue.scala 349:37:@44945.6]
  wire [31:0] _GEN_2270; // @[LoadQueue.scala 349:37:@44945.6]
  wire [31:0] _GEN_2271; // @[LoadQueue.scala 349:37:@44945.6]
  wire [31:0] _GEN_2272; // @[LoadQueue.scala 349:37:@44945.6]
  wire [31:0] _GEN_2273; // @[LoadQueue.scala 349:37:@44945.6]
  wire [31:0] _GEN_2274; // @[LoadQueue.scala 349:37:@44945.6]
  wire [31:0] _GEN_2275; // @[LoadQueue.scala 349:37:@44945.6]
  wire  _GEN_2279; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2280; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2281; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2282; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2283; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2284; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2285; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2286; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2287; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2288; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2289; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2290; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2291; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2292; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2293; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2295; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2296; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2297; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2298; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2299; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2300; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2301; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2302; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2303; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2304; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2305; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2306; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2307; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2308; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _GEN_2309; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _T_102167; // @[LoadQueue.scala 363:29:@44952.4]
  wire  _T_102168; // @[LoadQueue.scala 363:63:@44953.4]
  wire  _T_102170; // @[LoadQueue.scala 363:75:@44954.4]
  wire  _T_102171; // @[LoadQueue.scala 363:72:@44955.4]
  wire  _T_102172; // @[LoadQueue.scala 363:54:@44956.4]
  wire [4:0] _T_102175; // @[util.scala 10:8:@44958.6]
  wire [4:0] _GEN_544; // @[util.scala 10:14:@44959.6]
  wire [4:0] _T_102176; // @[util.scala 10:14:@44959.6]
  wire [4:0] _GEN_2310; // @[LoadQueue.scala 363:91:@44957.4]
  wire [3:0] _GEN_2408; // @[util.scala 10:8:@44963.6]
  wire [4:0] _T_102178; // @[util.scala 10:8:@44963.6]
  wire [4:0] _GEN_545; // @[util.scala 10:14:@44964.6]
  wire [4:0] _T_102179; // @[util.scala 10:14:@44964.6]
  wire [4:0] _GEN_2311; // @[LoadQueue.scala 367:20:@44962.4]
  wire  _T_102181; // @[LoadQueue.scala 371:82:@44967.4]
  wire  _T_102182; // @[LoadQueue.scala 371:79:@44968.4]
  wire  _T_102184; // @[LoadQueue.scala 371:82:@44969.4]
  wire  _T_102185; // @[LoadQueue.scala 371:79:@44970.4]
  wire  _T_102187; // @[LoadQueue.scala 371:82:@44971.4]
  wire  _T_102188; // @[LoadQueue.scala 371:79:@44972.4]
  wire  _T_102190; // @[LoadQueue.scala 371:82:@44973.4]
  wire  _T_102191; // @[LoadQueue.scala 371:79:@44974.4]
  wire  _T_102193; // @[LoadQueue.scala 371:82:@44975.4]
  wire  _T_102194; // @[LoadQueue.scala 371:79:@44976.4]
  wire  _T_102196; // @[LoadQueue.scala 371:82:@44977.4]
  wire  _T_102197; // @[LoadQueue.scala 371:79:@44978.4]
  wire  _T_102199; // @[LoadQueue.scala 371:82:@44979.4]
  wire  _T_102200; // @[LoadQueue.scala 371:79:@44980.4]
  wire  _T_102202; // @[LoadQueue.scala 371:82:@44981.4]
  wire  _T_102203; // @[LoadQueue.scala 371:79:@44982.4]
  wire  _T_102205; // @[LoadQueue.scala 371:82:@44983.4]
  wire  _T_102206; // @[LoadQueue.scala 371:79:@44984.4]
  wire  _T_102208; // @[LoadQueue.scala 371:82:@44985.4]
  wire  _T_102209; // @[LoadQueue.scala 371:79:@44986.4]
  wire  _T_102211; // @[LoadQueue.scala 371:82:@44987.4]
  wire  _T_102212; // @[LoadQueue.scala 371:79:@44988.4]
  wire  _T_102214; // @[LoadQueue.scala 371:82:@44989.4]
  wire  _T_102215; // @[LoadQueue.scala 371:79:@44990.4]
  wire  _T_102217; // @[LoadQueue.scala 371:82:@44991.4]
  wire  _T_102218; // @[LoadQueue.scala 371:79:@44992.4]
  wire  _T_102220; // @[LoadQueue.scala 371:82:@44993.4]
  wire  _T_102221; // @[LoadQueue.scala 371:79:@44994.4]
  wire  _T_102223; // @[LoadQueue.scala 371:82:@44995.4]
  wire  _T_102224; // @[LoadQueue.scala 371:79:@44996.4]
  wire  _T_102226; // @[LoadQueue.scala 371:82:@44997.4]
  wire  _T_102227; // @[LoadQueue.scala 371:79:@44998.4]
  wire  _T_102252; // @[LoadQueue.scala 371:96:@45017.4]
  wire  _T_102253; // @[LoadQueue.scala 371:96:@45018.4]
  wire  _T_102254; // @[LoadQueue.scala 371:96:@45019.4]
  wire  _T_102255; // @[LoadQueue.scala 371:96:@45020.4]
  wire  _T_102256; // @[LoadQueue.scala 371:96:@45021.4]
  wire  _T_102257; // @[LoadQueue.scala 371:96:@45022.4]
  wire  _T_102258; // @[LoadQueue.scala 371:96:@45023.4]
  wire  _T_102259; // @[LoadQueue.scala 371:96:@45024.4]
  wire  _T_102260; // @[LoadQueue.scala 371:96:@45025.4]
  wire  _T_102261; // @[LoadQueue.scala 371:96:@45026.4]
  wire  _T_102262; // @[LoadQueue.scala 371:96:@45027.4]
  wire  _T_102263; // @[LoadQueue.scala 371:96:@45028.4]
  wire  _T_102264; // @[LoadQueue.scala 371:96:@45029.4]
  wire  _T_102265; // @[LoadQueue.scala 371:96:@45030.4]
  assign _GEN_2312 = {{2'd0}, tail}; // @[util.scala 14:20:@5032.4]
  assign _T_1724 = 6'h10 - _GEN_2312; // @[util.scala 14:20:@5032.4]
  assign _T_1725 = $unsigned(_T_1724); // @[util.scala 14:20:@5033.4]
  assign _T_1726 = _T_1725[5:0]; // @[util.scala 14:20:@5034.4]
  assign _GEN_0 = _T_1726 % 6'h10; // @[util.scala 14:25:@5035.4]
  assign _T_1727 = _GEN_0[4:0]; // @[util.scala 14:25:@5035.4]
  assign _GEN_2313 = {{3'd0}, io_bbNumLoads}; // @[LoadQueue.scala 71:46:@5036.4]
  assign _T_1728 = _T_1727 < _GEN_2313; // @[LoadQueue.scala 71:46:@5036.4]
  assign initBits_0 = _T_1728 & io_bbStart; // @[LoadQueue.scala 71:63:@5037.4]
  assign _T_1733 = 6'h11 - _GEN_2312; // @[util.scala 14:20:@5039.4]
  assign _T_1734 = $unsigned(_T_1733); // @[util.scala 14:20:@5040.4]
  assign _T_1735 = _T_1734[5:0]; // @[util.scala 14:20:@5041.4]
  assign _GEN_16 = _T_1735 % 6'h10; // @[util.scala 14:25:@5042.4]
  assign _T_1736 = _GEN_16[4:0]; // @[util.scala 14:25:@5042.4]
  assign _T_1737 = _T_1736 < _GEN_2313; // @[LoadQueue.scala 71:46:@5043.4]
  assign initBits_1 = _T_1737 & io_bbStart; // @[LoadQueue.scala 71:63:@5044.4]
  assign _T_1742 = 6'h12 - _GEN_2312; // @[util.scala 14:20:@5046.4]
  assign _T_1743 = $unsigned(_T_1742); // @[util.scala 14:20:@5047.4]
  assign _T_1744 = _T_1743[5:0]; // @[util.scala 14:20:@5048.4]
  assign _GEN_34 = _T_1744 % 6'h10; // @[util.scala 14:25:@5049.4]
  assign _T_1745 = _GEN_34[4:0]; // @[util.scala 14:25:@5049.4]
  assign _T_1746 = _T_1745 < _GEN_2313; // @[LoadQueue.scala 71:46:@5050.4]
  assign initBits_2 = _T_1746 & io_bbStart; // @[LoadQueue.scala 71:63:@5051.4]
  assign _T_1751 = 6'h13 - _GEN_2312; // @[util.scala 14:20:@5053.4]
  assign _T_1752 = $unsigned(_T_1751); // @[util.scala 14:20:@5054.4]
  assign _T_1753 = _T_1752[5:0]; // @[util.scala 14:20:@5055.4]
  assign _GEN_50 = _T_1753 % 6'h10; // @[util.scala 14:25:@5056.4]
  assign _T_1754 = _GEN_50[4:0]; // @[util.scala 14:25:@5056.4]
  assign _T_1755 = _T_1754 < _GEN_2313; // @[LoadQueue.scala 71:46:@5057.4]
  assign initBits_3 = _T_1755 & io_bbStart; // @[LoadQueue.scala 71:63:@5058.4]
  assign _T_1760 = 6'h14 - _GEN_2312; // @[util.scala 14:20:@5060.4]
  assign _T_1761 = $unsigned(_T_1760); // @[util.scala 14:20:@5061.4]
  assign _T_1762 = _T_1761[5:0]; // @[util.scala 14:20:@5062.4]
  assign _GEN_68 = _T_1762 % 6'h10; // @[util.scala 14:25:@5063.4]
  assign _T_1763 = _GEN_68[4:0]; // @[util.scala 14:25:@5063.4]
  assign _T_1764 = _T_1763 < _GEN_2313; // @[LoadQueue.scala 71:46:@5064.4]
  assign initBits_4 = _T_1764 & io_bbStart; // @[LoadQueue.scala 71:63:@5065.4]
  assign _T_1769 = 6'h15 - _GEN_2312; // @[util.scala 14:20:@5067.4]
  assign _T_1770 = $unsigned(_T_1769); // @[util.scala 14:20:@5068.4]
  assign _T_1771 = _T_1770[5:0]; // @[util.scala 14:20:@5069.4]
  assign _GEN_84 = _T_1771 % 6'h10; // @[util.scala 14:25:@5070.4]
  assign _T_1772 = _GEN_84[4:0]; // @[util.scala 14:25:@5070.4]
  assign _T_1773 = _T_1772 < _GEN_2313; // @[LoadQueue.scala 71:46:@5071.4]
  assign initBits_5 = _T_1773 & io_bbStart; // @[LoadQueue.scala 71:63:@5072.4]
  assign _T_1778 = 6'h16 - _GEN_2312; // @[util.scala 14:20:@5074.4]
  assign _T_1779 = $unsigned(_T_1778); // @[util.scala 14:20:@5075.4]
  assign _T_1780 = _T_1779[5:0]; // @[util.scala 14:20:@5076.4]
  assign _GEN_102 = _T_1780 % 6'h10; // @[util.scala 14:25:@5077.4]
  assign _T_1781 = _GEN_102[4:0]; // @[util.scala 14:25:@5077.4]
  assign _T_1782 = _T_1781 < _GEN_2313; // @[LoadQueue.scala 71:46:@5078.4]
  assign initBits_6 = _T_1782 & io_bbStart; // @[LoadQueue.scala 71:63:@5079.4]
  assign _T_1787 = 6'h17 - _GEN_2312; // @[util.scala 14:20:@5081.4]
  assign _T_1788 = $unsigned(_T_1787); // @[util.scala 14:20:@5082.4]
  assign _T_1789 = _T_1788[5:0]; // @[util.scala 14:20:@5083.4]
  assign _GEN_118 = _T_1789 % 6'h10; // @[util.scala 14:25:@5084.4]
  assign _T_1790 = _GEN_118[4:0]; // @[util.scala 14:25:@5084.4]
  assign _T_1791 = _T_1790 < _GEN_2313; // @[LoadQueue.scala 71:46:@5085.4]
  assign initBits_7 = _T_1791 & io_bbStart; // @[LoadQueue.scala 71:63:@5086.4]
  assign _T_1796 = 6'h18 - _GEN_2312; // @[util.scala 14:20:@5088.4]
  assign _T_1797 = $unsigned(_T_1796); // @[util.scala 14:20:@5089.4]
  assign _T_1798 = _T_1797[5:0]; // @[util.scala 14:20:@5090.4]
  assign _GEN_136 = _T_1798 % 6'h10; // @[util.scala 14:25:@5091.4]
  assign _T_1799 = _GEN_136[4:0]; // @[util.scala 14:25:@5091.4]
  assign _T_1800 = _T_1799 < _GEN_2313; // @[LoadQueue.scala 71:46:@5092.4]
  assign initBits_8 = _T_1800 & io_bbStart; // @[LoadQueue.scala 71:63:@5093.4]
  assign _T_1805 = 6'h19 - _GEN_2312; // @[util.scala 14:20:@5095.4]
  assign _T_1806 = $unsigned(_T_1805); // @[util.scala 14:20:@5096.4]
  assign _T_1807 = _T_1806[5:0]; // @[util.scala 14:20:@5097.4]
  assign _GEN_152 = _T_1807 % 6'h10; // @[util.scala 14:25:@5098.4]
  assign _T_1808 = _GEN_152[4:0]; // @[util.scala 14:25:@5098.4]
  assign _T_1809 = _T_1808 < _GEN_2313; // @[LoadQueue.scala 71:46:@5099.4]
  assign initBits_9 = _T_1809 & io_bbStart; // @[LoadQueue.scala 71:63:@5100.4]
  assign _T_1814 = 6'h1a - _GEN_2312; // @[util.scala 14:20:@5102.4]
  assign _T_1815 = $unsigned(_T_1814); // @[util.scala 14:20:@5103.4]
  assign _T_1816 = _T_1815[5:0]; // @[util.scala 14:20:@5104.4]
  assign _GEN_170 = _T_1816 % 6'h10; // @[util.scala 14:25:@5105.4]
  assign _T_1817 = _GEN_170[4:0]; // @[util.scala 14:25:@5105.4]
  assign _T_1818 = _T_1817 < _GEN_2313; // @[LoadQueue.scala 71:46:@5106.4]
  assign initBits_10 = _T_1818 & io_bbStart; // @[LoadQueue.scala 71:63:@5107.4]
  assign _T_1823 = 6'h1b - _GEN_2312; // @[util.scala 14:20:@5109.4]
  assign _T_1824 = $unsigned(_T_1823); // @[util.scala 14:20:@5110.4]
  assign _T_1825 = _T_1824[5:0]; // @[util.scala 14:20:@5111.4]
  assign _GEN_186 = _T_1825 % 6'h10; // @[util.scala 14:25:@5112.4]
  assign _T_1826 = _GEN_186[4:0]; // @[util.scala 14:25:@5112.4]
  assign _T_1827 = _T_1826 < _GEN_2313; // @[LoadQueue.scala 71:46:@5113.4]
  assign initBits_11 = _T_1827 & io_bbStart; // @[LoadQueue.scala 71:63:@5114.4]
  assign _T_1832 = 6'h1c - _GEN_2312; // @[util.scala 14:20:@5116.4]
  assign _T_1833 = $unsigned(_T_1832); // @[util.scala 14:20:@5117.4]
  assign _T_1834 = _T_1833[5:0]; // @[util.scala 14:20:@5118.4]
  assign _GEN_204 = _T_1834 % 6'h10; // @[util.scala 14:25:@5119.4]
  assign _T_1835 = _GEN_204[4:0]; // @[util.scala 14:25:@5119.4]
  assign _T_1836 = _T_1835 < _GEN_2313; // @[LoadQueue.scala 71:46:@5120.4]
  assign initBits_12 = _T_1836 & io_bbStart; // @[LoadQueue.scala 71:63:@5121.4]
  assign _T_1841 = 6'h1d - _GEN_2312; // @[util.scala 14:20:@5123.4]
  assign _T_1842 = $unsigned(_T_1841); // @[util.scala 14:20:@5124.4]
  assign _T_1843 = _T_1842[5:0]; // @[util.scala 14:20:@5125.4]
  assign _GEN_220 = _T_1843 % 6'h10; // @[util.scala 14:25:@5126.4]
  assign _T_1844 = _GEN_220[4:0]; // @[util.scala 14:25:@5126.4]
  assign _T_1845 = _T_1844 < _GEN_2313; // @[LoadQueue.scala 71:46:@5127.4]
  assign initBits_13 = _T_1845 & io_bbStart; // @[LoadQueue.scala 71:63:@5128.4]
  assign _T_1850 = 6'h1e - _GEN_2312; // @[util.scala 14:20:@5130.4]
  assign _T_1851 = $unsigned(_T_1850); // @[util.scala 14:20:@5131.4]
  assign _T_1852 = _T_1851[5:0]; // @[util.scala 14:20:@5132.4]
  assign _GEN_238 = _T_1852 % 6'h10; // @[util.scala 14:25:@5133.4]
  assign _T_1853 = _GEN_238[4:0]; // @[util.scala 14:25:@5133.4]
  assign _T_1854 = _T_1853 < _GEN_2313; // @[LoadQueue.scala 71:46:@5134.4]
  assign initBits_14 = _T_1854 & io_bbStart; // @[LoadQueue.scala 71:63:@5135.4]
  assign _T_1859 = 6'h1f - _GEN_2312; // @[util.scala 14:20:@5137.4]
  assign _T_1860 = $unsigned(_T_1859); // @[util.scala 14:20:@5138.4]
  assign _T_1861 = _T_1860[5:0]; // @[util.scala 14:20:@5139.4]
  assign _GEN_254 = _T_1861 % 6'h10; // @[util.scala 14:25:@5140.4]
  assign _T_1862 = _GEN_254[4:0]; // @[util.scala 14:25:@5140.4]
  assign _T_1863 = _T_1862 < _GEN_2313; // @[LoadQueue.scala 71:46:@5141.4]
  assign initBits_15 = _T_1863 & io_bbStart; // @[LoadQueue.scala 71:63:@5142.4]
  assign _T_1886 = allocatedEntries_0 | initBits_0; // @[LoadQueue.scala 73:78:@5160.4]
  assign _T_1887 = allocatedEntries_1 | initBits_1; // @[LoadQueue.scala 73:78:@5161.4]
  assign _T_1888 = allocatedEntries_2 | initBits_2; // @[LoadQueue.scala 73:78:@5162.4]
  assign _T_1889 = allocatedEntries_3 | initBits_3; // @[LoadQueue.scala 73:78:@5163.4]
  assign _T_1890 = allocatedEntries_4 | initBits_4; // @[LoadQueue.scala 73:78:@5164.4]
  assign _T_1891 = allocatedEntries_5 | initBits_5; // @[LoadQueue.scala 73:78:@5165.4]
  assign _T_1892 = allocatedEntries_6 | initBits_6; // @[LoadQueue.scala 73:78:@5166.4]
  assign _T_1893 = allocatedEntries_7 | initBits_7; // @[LoadQueue.scala 73:78:@5167.4]
  assign _T_1894 = allocatedEntries_8 | initBits_8; // @[LoadQueue.scala 73:78:@5168.4]
  assign _T_1895 = allocatedEntries_9 | initBits_9; // @[LoadQueue.scala 73:78:@5169.4]
  assign _T_1896 = allocatedEntries_10 | initBits_10; // @[LoadQueue.scala 73:78:@5170.4]
  assign _T_1897 = allocatedEntries_11 | initBits_11; // @[LoadQueue.scala 73:78:@5171.4]
  assign _T_1898 = allocatedEntries_12 | initBits_12; // @[LoadQueue.scala 73:78:@5172.4]
  assign _T_1899 = allocatedEntries_13 | initBits_13; // @[LoadQueue.scala 73:78:@5173.4]
  assign _T_1900 = allocatedEntries_14 | initBits_14; // @[LoadQueue.scala 73:78:@5174.4]
  assign _T_1901 = allocatedEntries_15 | initBits_15; // @[LoadQueue.scala 73:78:@5175.4]
  assign _T_1932 = _T_1727[3:0]; // @[:@5215.6]
  assign _GEN_1 = 4'h1 == _T_1932 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_2 = 4'h2 == _T_1932 ? io_bbLoadOffsets_2 : _GEN_1; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_3 = 4'h3 == _T_1932 ? io_bbLoadOffsets_3 : _GEN_2; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_4 = 4'h4 == _T_1932 ? io_bbLoadOffsets_4 : _GEN_3; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_5 = 4'h5 == _T_1932 ? io_bbLoadOffsets_5 : _GEN_4; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_6 = 4'h6 == _T_1932 ? io_bbLoadOffsets_6 : _GEN_5; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_7 = 4'h7 == _T_1932 ? io_bbLoadOffsets_7 : _GEN_6; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_8 = 4'h8 == _T_1932 ? io_bbLoadOffsets_8 : _GEN_7; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_9 = 4'h9 == _T_1932 ? io_bbLoadOffsets_9 : _GEN_8; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_10 = 4'ha == _T_1932 ? io_bbLoadOffsets_10 : _GEN_9; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_11 = 4'hb == _T_1932 ? io_bbLoadOffsets_11 : _GEN_10; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_12 = 4'hc == _T_1932 ? io_bbLoadOffsets_12 : _GEN_11; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_13 = 4'hd == _T_1932 ? io_bbLoadOffsets_13 : _GEN_12; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_14 = 4'he == _T_1932 ? io_bbLoadOffsets_14 : _GEN_13; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_15 = 4'hf == _T_1932 ? io_bbLoadOffsets_15 : _GEN_14; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_17 = 4'h1 == _T_1932 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@5223.6]
  assign _GEN_18 = 4'h2 == _T_1932 ? 1'h0 : _GEN_17; // @[LoadQueue.scala 78:18:@5223.6]
  assign _GEN_19 = 4'h3 == _T_1932 ? 1'h0 : _GEN_18; // @[LoadQueue.scala 78:18:@5223.6]
  assign _GEN_20 = 4'h4 == _T_1932 ? 1'h0 : _GEN_19; // @[LoadQueue.scala 78:18:@5223.6]
  assign _GEN_21 = 4'h5 == _T_1932 ? 1'h0 : _GEN_20; // @[LoadQueue.scala 78:18:@5223.6]
  assign _GEN_22 = 4'h6 == _T_1932 ? 1'h0 : _GEN_21; // @[LoadQueue.scala 78:18:@5223.6]
  assign _GEN_23 = 4'h7 == _T_1932 ? 1'h0 : _GEN_22; // @[LoadQueue.scala 78:18:@5223.6]
  assign _GEN_24 = 4'h8 == _T_1932 ? 1'h0 : _GEN_23; // @[LoadQueue.scala 78:18:@5223.6]
  assign _GEN_25 = 4'h9 == _T_1932 ? 1'h0 : _GEN_24; // @[LoadQueue.scala 78:18:@5223.6]
  assign _GEN_26 = 4'ha == _T_1932 ? 1'h0 : _GEN_25; // @[LoadQueue.scala 78:18:@5223.6]
  assign _GEN_27 = 4'hb == _T_1932 ? 1'h0 : _GEN_26; // @[LoadQueue.scala 78:18:@5223.6]
  assign _GEN_28 = 4'hc == _T_1932 ? 1'h0 : _GEN_27; // @[LoadQueue.scala 78:18:@5223.6]
  assign _GEN_29 = 4'hd == _T_1932 ? 1'h0 : _GEN_28; // @[LoadQueue.scala 78:18:@5223.6]
  assign _GEN_30 = 4'he == _T_1932 ? 1'h0 : _GEN_29; // @[LoadQueue.scala 78:18:@5223.6]
  assign _GEN_31 = 4'hf == _T_1932 ? 1'h0 : _GEN_30; // @[LoadQueue.scala 78:18:@5223.6]
  assign _GEN_32 = initBits_0 ? _GEN_15 : offsetQ_0; // @[LoadQueue.scala 76:25:@5209.4]
  assign _GEN_33 = initBits_0 ? _GEN_31 : portQ_0; // @[LoadQueue.scala 76:25:@5209.4]
  assign _T_1950 = _T_1736[3:0]; // @[:@5231.6]
  assign _GEN_35 = 4'h1 == _T_1950 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_36 = 4'h2 == _T_1950 ? io_bbLoadOffsets_2 : _GEN_35; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_37 = 4'h3 == _T_1950 ? io_bbLoadOffsets_3 : _GEN_36; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_38 = 4'h4 == _T_1950 ? io_bbLoadOffsets_4 : _GEN_37; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_39 = 4'h5 == _T_1950 ? io_bbLoadOffsets_5 : _GEN_38; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_40 = 4'h6 == _T_1950 ? io_bbLoadOffsets_6 : _GEN_39; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_41 = 4'h7 == _T_1950 ? io_bbLoadOffsets_7 : _GEN_40; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_42 = 4'h8 == _T_1950 ? io_bbLoadOffsets_8 : _GEN_41; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_43 = 4'h9 == _T_1950 ? io_bbLoadOffsets_9 : _GEN_42; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_44 = 4'ha == _T_1950 ? io_bbLoadOffsets_10 : _GEN_43; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_45 = 4'hb == _T_1950 ? io_bbLoadOffsets_11 : _GEN_44; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_46 = 4'hc == _T_1950 ? io_bbLoadOffsets_12 : _GEN_45; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_47 = 4'hd == _T_1950 ? io_bbLoadOffsets_13 : _GEN_46; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_48 = 4'he == _T_1950 ? io_bbLoadOffsets_14 : _GEN_47; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_49 = 4'hf == _T_1950 ? io_bbLoadOffsets_15 : _GEN_48; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_51 = 4'h1 == _T_1950 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@5239.6]
  assign _GEN_52 = 4'h2 == _T_1950 ? 1'h0 : _GEN_51; // @[LoadQueue.scala 78:18:@5239.6]
  assign _GEN_53 = 4'h3 == _T_1950 ? 1'h0 : _GEN_52; // @[LoadQueue.scala 78:18:@5239.6]
  assign _GEN_54 = 4'h4 == _T_1950 ? 1'h0 : _GEN_53; // @[LoadQueue.scala 78:18:@5239.6]
  assign _GEN_55 = 4'h5 == _T_1950 ? 1'h0 : _GEN_54; // @[LoadQueue.scala 78:18:@5239.6]
  assign _GEN_56 = 4'h6 == _T_1950 ? 1'h0 : _GEN_55; // @[LoadQueue.scala 78:18:@5239.6]
  assign _GEN_57 = 4'h7 == _T_1950 ? 1'h0 : _GEN_56; // @[LoadQueue.scala 78:18:@5239.6]
  assign _GEN_58 = 4'h8 == _T_1950 ? 1'h0 : _GEN_57; // @[LoadQueue.scala 78:18:@5239.6]
  assign _GEN_59 = 4'h9 == _T_1950 ? 1'h0 : _GEN_58; // @[LoadQueue.scala 78:18:@5239.6]
  assign _GEN_60 = 4'ha == _T_1950 ? 1'h0 : _GEN_59; // @[LoadQueue.scala 78:18:@5239.6]
  assign _GEN_61 = 4'hb == _T_1950 ? 1'h0 : _GEN_60; // @[LoadQueue.scala 78:18:@5239.6]
  assign _GEN_62 = 4'hc == _T_1950 ? 1'h0 : _GEN_61; // @[LoadQueue.scala 78:18:@5239.6]
  assign _GEN_63 = 4'hd == _T_1950 ? 1'h0 : _GEN_62; // @[LoadQueue.scala 78:18:@5239.6]
  assign _GEN_64 = 4'he == _T_1950 ? 1'h0 : _GEN_63; // @[LoadQueue.scala 78:18:@5239.6]
  assign _GEN_65 = 4'hf == _T_1950 ? 1'h0 : _GEN_64; // @[LoadQueue.scala 78:18:@5239.6]
  assign _GEN_66 = initBits_1 ? _GEN_49 : offsetQ_1; // @[LoadQueue.scala 76:25:@5225.4]
  assign _GEN_67 = initBits_1 ? _GEN_65 : portQ_1; // @[LoadQueue.scala 76:25:@5225.4]
  assign _T_1968 = _T_1745[3:0]; // @[:@5247.6]
  assign _GEN_69 = 4'h1 == _T_1968 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_70 = 4'h2 == _T_1968 ? io_bbLoadOffsets_2 : _GEN_69; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_71 = 4'h3 == _T_1968 ? io_bbLoadOffsets_3 : _GEN_70; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_72 = 4'h4 == _T_1968 ? io_bbLoadOffsets_4 : _GEN_71; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_73 = 4'h5 == _T_1968 ? io_bbLoadOffsets_5 : _GEN_72; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_74 = 4'h6 == _T_1968 ? io_bbLoadOffsets_6 : _GEN_73; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_75 = 4'h7 == _T_1968 ? io_bbLoadOffsets_7 : _GEN_74; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_76 = 4'h8 == _T_1968 ? io_bbLoadOffsets_8 : _GEN_75; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_77 = 4'h9 == _T_1968 ? io_bbLoadOffsets_9 : _GEN_76; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_78 = 4'ha == _T_1968 ? io_bbLoadOffsets_10 : _GEN_77; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_79 = 4'hb == _T_1968 ? io_bbLoadOffsets_11 : _GEN_78; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_80 = 4'hc == _T_1968 ? io_bbLoadOffsets_12 : _GEN_79; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_81 = 4'hd == _T_1968 ? io_bbLoadOffsets_13 : _GEN_80; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_82 = 4'he == _T_1968 ? io_bbLoadOffsets_14 : _GEN_81; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_83 = 4'hf == _T_1968 ? io_bbLoadOffsets_15 : _GEN_82; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_85 = 4'h1 == _T_1968 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@5255.6]
  assign _GEN_86 = 4'h2 == _T_1968 ? 1'h0 : _GEN_85; // @[LoadQueue.scala 78:18:@5255.6]
  assign _GEN_87 = 4'h3 == _T_1968 ? 1'h0 : _GEN_86; // @[LoadQueue.scala 78:18:@5255.6]
  assign _GEN_88 = 4'h4 == _T_1968 ? 1'h0 : _GEN_87; // @[LoadQueue.scala 78:18:@5255.6]
  assign _GEN_89 = 4'h5 == _T_1968 ? 1'h0 : _GEN_88; // @[LoadQueue.scala 78:18:@5255.6]
  assign _GEN_90 = 4'h6 == _T_1968 ? 1'h0 : _GEN_89; // @[LoadQueue.scala 78:18:@5255.6]
  assign _GEN_91 = 4'h7 == _T_1968 ? 1'h0 : _GEN_90; // @[LoadQueue.scala 78:18:@5255.6]
  assign _GEN_92 = 4'h8 == _T_1968 ? 1'h0 : _GEN_91; // @[LoadQueue.scala 78:18:@5255.6]
  assign _GEN_93 = 4'h9 == _T_1968 ? 1'h0 : _GEN_92; // @[LoadQueue.scala 78:18:@5255.6]
  assign _GEN_94 = 4'ha == _T_1968 ? 1'h0 : _GEN_93; // @[LoadQueue.scala 78:18:@5255.6]
  assign _GEN_95 = 4'hb == _T_1968 ? 1'h0 : _GEN_94; // @[LoadQueue.scala 78:18:@5255.6]
  assign _GEN_96 = 4'hc == _T_1968 ? 1'h0 : _GEN_95; // @[LoadQueue.scala 78:18:@5255.6]
  assign _GEN_97 = 4'hd == _T_1968 ? 1'h0 : _GEN_96; // @[LoadQueue.scala 78:18:@5255.6]
  assign _GEN_98 = 4'he == _T_1968 ? 1'h0 : _GEN_97; // @[LoadQueue.scala 78:18:@5255.6]
  assign _GEN_99 = 4'hf == _T_1968 ? 1'h0 : _GEN_98; // @[LoadQueue.scala 78:18:@5255.6]
  assign _GEN_100 = initBits_2 ? _GEN_83 : offsetQ_2; // @[LoadQueue.scala 76:25:@5241.4]
  assign _GEN_101 = initBits_2 ? _GEN_99 : portQ_2; // @[LoadQueue.scala 76:25:@5241.4]
  assign _T_1986 = _T_1754[3:0]; // @[:@5263.6]
  assign _GEN_103 = 4'h1 == _T_1986 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_104 = 4'h2 == _T_1986 ? io_bbLoadOffsets_2 : _GEN_103; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_105 = 4'h3 == _T_1986 ? io_bbLoadOffsets_3 : _GEN_104; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_106 = 4'h4 == _T_1986 ? io_bbLoadOffsets_4 : _GEN_105; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_107 = 4'h5 == _T_1986 ? io_bbLoadOffsets_5 : _GEN_106; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_108 = 4'h6 == _T_1986 ? io_bbLoadOffsets_6 : _GEN_107; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_109 = 4'h7 == _T_1986 ? io_bbLoadOffsets_7 : _GEN_108; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_110 = 4'h8 == _T_1986 ? io_bbLoadOffsets_8 : _GEN_109; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_111 = 4'h9 == _T_1986 ? io_bbLoadOffsets_9 : _GEN_110; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_112 = 4'ha == _T_1986 ? io_bbLoadOffsets_10 : _GEN_111; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_113 = 4'hb == _T_1986 ? io_bbLoadOffsets_11 : _GEN_112; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_114 = 4'hc == _T_1986 ? io_bbLoadOffsets_12 : _GEN_113; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_115 = 4'hd == _T_1986 ? io_bbLoadOffsets_13 : _GEN_114; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_116 = 4'he == _T_1986 ? io_bbLoadOffsets_14 : _GEN_115; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_117 = 4'hf == _T_1986 ? io_bbLoadOffsets_15 : _GEN_116; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_119 = 4'h1 == _T_1986 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@5271.6]
  assign _GEN_120 = 4'h2 == _T_1986 ? 1'h0 : _GEN_119; // @[LoadQueue.scala 78:18:@5271.6]
  assign _GEN_121 = 4'h3 == _T_1986 ? 1'h0 : _GEN_120; // @[LoadQueue.scala 78:18:@5271.6]
  assign _GEN_122 = 4'h4 == _T_1986 ? 1'h0 : _GEN_121; // @[LoadQueue.scala 78:18:@5271.6]
  assign _GEN_123 = 4'h5 == _T_1986 ? 1'h0 : _GEN_122; // @[LoadQueue.scala 78:18:@5271.6]
  assign _GEN_124 = 4'h6 == _T_1986 ? 1'h0 : _GEN_123; // @[LoadQueue.scala 78:18:@5271.6]
  assign _GEN_125 = 4'h7 == _T_1986 ? 1'h0 : _GEN_124; // @[LoadQueue.scala 78:18:@5271.6]
  assign _GEN_126 = 4'h8 == _T_1986 ? 1'h0 : _GEN_125; // @[LoadQueue.scala 78:18:@5271.6]
  assign _GEN_127 = 4'h9 == _T_1986 ? 1'h0 : _GEN_126; // @[LoadQueue.scala 78:18:@5271.6]
  assign _GEN_128 = 4'ha == _T_1986 ? 1'h0 : _GEN_127; // @[LoadQueue.scala 78:18:@5271.6]
  assign _GEN_129 = 4'hb == _T_1986 ? 1'h0 : _GEN_128; // @[LoadQueue.scala 78:18:@5271.6]
  assign _GEN_130 = 4'hc == _T_1986 ? 1'h0 : _GEN_129; // @[LoadQueue.scala 78:18:@5271.6]
  assign _GEN_131 = 4'hd == _T_1986 ? 1'h0 : _GEN_130; // @[LoadQueue.scala 78:18:@5271.6]
  assign _GEN_132 = 4'he == _T_1986 ? 1'h0 : _GEN_131; // @[LoadQueue.scala 78:18:@5271.6]
  assign _GEN_133 = 4'hf == _T_1986 ? 1'h0 : _GEN_132; // @[LoadQueue.scala 78:18:@5271.6]
  assign _GEN_134 = initBits_3 ? _GEN_117 : offsetQ_3; // @[LoadQueue.scala 76:25:@5257.4]
  assign _GEN_135 = initBits_3 ? _GEN_133 : portQ_3; // @[LoadQueue.scala 76:25:@5257.4]
  assign _T_2004 = _T_1763[3:0]; // @[:@5279.6]
  assign _GEN_137 = 4'h1 == _T_2004 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_138 = 4'h2 == _T_2004 ? io_bbLoadOffsets_2 : _GEN_137; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_139 = 4'h3 == _T_2004 ? io_bbLoadOffsets_3 : _GEN_138; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_140 = 4'h4 == _T_2004 ? io_bbLoadOffsets_4 : _GEN_139; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_141 = 4'h5 == _T_2004 ? io_bbLoadOffsets_5 : _GEN_140; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_142 = 4'h6 == _T_2004 ? io_bbLoadOffsets_6 : _GEN_141; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_143 = 4'h7 == _T_2004 ? io_bbLoadOffsets_7 : _GEN_142; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_144 = 4'h8 == _T_2004 ? io_bbLoadOffsets_8 : _GEN_143; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_145 = 4'h9 == _T_2004 ? io_bbLoadOffsets_9 : _GEN_144; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_146 = 4'ha == _T_2004 ? io_bbLoadOffsets_10 : _GEN_145; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_147 = 4'hb == _T_2004 ? io_bbLoadOffsets_11 : _GEN_146; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_148 = 4'hc == _T_2004 ? io_bbLoadOffsets_12 : _GEN_147; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_149 = 4'hd == _T_2004 ? io_bbLoadOffsets_13 : _GEN_148; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_150 = 4'he == _T_2004 ? io_bbLoadOffsets_14 : _GEN_149; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_151 = 4'hf == _T_2004 ? io_bbLoadOffsets_15 : _GEN_150; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_153 = 4'h1 == _T_2004 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@5287.6]
  assign _GEN_154 = 4'h2 == _T_2004 ? 1'h0 : _GEN_153; // @[LoadQueue.scala 78:18:@5287.6]
  assign _GEN_155 = 4'h3 == _T_2004 ? 1'h0 : _GEN_154; // @[LoadQueue.scala 78:18:@5287.6]
  assign _GEN_156 = 4'h4 == _T_2004 ? 1'h0 : _GEN_155; // @[LoadQueue.scala 78:18:@5287.6]
  assign _GEN_157 = 4'h5 == _T_2004 ? 1'h0 : _GEN_156; // @[LoadQueue.scala 78:18:@5287.6]
  assign _GEN_158 = 4'h6 == _T_2004 ? 1'h0 : _GEN_157; // @[LoadQueue.scala 78:18:@5287.6]
  assign _GEN_159 = 4'h7 == _T_2004 ? 1'h0 : _GEN_158; // @[LoadQueue.scala 78:18:@5287.6]
  assign _GEN_160 = 4'h8 == _T_2004 ? 1'h0 : _GEN_159; // @[LoadQueue.scala 78:18:@5287.6]
  assign _GEN_161 = 4'h9 == _T_2004 ? 1'h0 : _GEN_160; // @[LoadQueue.scala 78:18:@5287.6]
  assign _GEN_162 = 4'ha == _T_2004 ? 1'h0 : _GEN_161; // @[LoadQueue.scala 78:18:@5287.6]
  assign _GEN_163 = 4'hb == _T_2004 ? 1'h0 : _GEN_162; // @[LoadQueue.scala 78:18:@5287.6]
  assign _GEN_164 = 4'hc == _T_2004 ? 1'h0 : _GEN_163; // @[LoadQueue.scala 78:18:@5287.6]
  assign _GEN_165 = 4'hd == _T_2004 ? 1'h0 : _GEN_164; // @[LoadQueue.scala 78:18:@5287.6]
  assign _GEN_166 = 4'he == _T_2004 ? 1'h0 : _GEN_165; // @[LoadQueue.scala 78:18:@5287.6]
  assign _GEN_167 = 4'hf == _T_2004 ? 1'h0 : _GEN_166; // @[LoadQueue.scala 78:18:@5287.6]
  assign _GEN_168 = initBits_4 ? _GEN_151 : offsetQ_4; // @[LoadQueue.scala 76:25:@5273.4]
  assign _GEN_169 = initBits_4 ? _GEN_167 : portQ_4; // @[LoadQueue.scala 76:25:@5273.4]
  assign _T_2022 = _T_1772[3:0]; // @[:@5295.6]
  assign _GEN_171 = 4'h1 == _T_2022 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_172 = 4'h2 == _T_2022 ? io_bbLoadOffsets_2 : _GEN_171; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_173 = 4'h3 == _T_2022 ? io_bbLoadOffsets_3 : _GEN_172; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_174 = 4'h4 == _T_2022 ? io_bbLoadOffsets_4 : _GEN_173; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_175 = 4'h5 == _T_2022 ? io_bbLoadOffsets_5 : _GEN_174; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_176 = 4'h6 == _T_2022 ? io_bbLoadOffsets_6 : _GEN_175; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_177 = 4'h7 == _T_2022 ? io_bbLoadOffsets_7 : _GEN_176; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_178 = 4'h8 == _T_2022 ? io_bbLoadOffsets_8 : _GEN_177; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_179 = 4'h9 == _T_2022 ? io_bbLoadOffsets_9 : _GEN_178; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_180 = 4'ha == _T_2022 ? io_bbLoadOffsets_10 : _GEN_179; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_181 = 4'hb == _T_2022 ? io_bbLoadOffsets_11 : _GEN_180; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_182 = 4'hc == _T_2022 ? io_bbLoadOffsets_12 : _GEN_181; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_183 = 4'hd == _T_2022 ? io_bbLoadOffsets_13 : _GEN_182; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_184 = 4'he == _T_2022 ? io_bbLoadOffsets_14 : _GEN_183; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_185 = 4'hf == _T_2022 ? io_bbLoadOffsets_15 : _GEN_184; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_187 = 4'h1 == _T_2022 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@5303.6]
  assign _GEN_188 = 4'h2 == _T_2022 ? 1'h0 : _GEN_187; // @[LoadQueue.scala 78:18:@5303.6]
  assign _GEN_189 = 4'h3 == _T_2022 ? 1'h0 : _GEN_188; // @[LoadQueue.scala 78:18:@5303.6]
  assign _GEN_190 = 4'h4 == _T_2022 ? 1'h0 : _GEN_189; // @[LoadQueue.scala 78:18:@5303.6]
  assign _GEN_191 = 4'h5 == _T_2022 ? 1'h0 : _GEN_190; // @[LoadQueue.scala 78:18:@5303.6]
  assign _GEN_192 = 4'h6 == _T_2022 ? 1'h0 : _GEN_191; // @[LoadQueue.scala 78:18:@5303.6]
  assign _GEN_193 = 4'h7 == _T_2022 ? 1'h0 : _GEN_192; // @[LoadQueue.scala 78:18:@5303.6]
  assign _GEN_194 = 4'h8 == _T_2022 ? 1'h0 : _GEN_193; // @[LoadQueue.scala 78:18:@5303.6]
  assign _GEN_195 = 4'h9 == _T_2022 ? 1'h0 : _GEN_194; // @[LoadQueue.scala 78:18:@5303.6]
  assign _GEN_196 = 4'ha == _T_2022 ? 1'h0 : _GEN_195; // @[LoadQueue.scala 78:18:@5303.6]
  assign _GEN_197 = 4'hb == _T_2022 ? 1'h0 : _GEN_196; // @[LoadQueue.scala 78:18:@5303.6]
  assign _GEN_198 = 4'hc == _T_2022 ? 1'h0 : _GEN_197; // @[LoadQueue.scala 78:18:@5303.6]
  assign _GEN_199 = 4'hd == _T_2022 ? 1'h0 : _GEN_198; // @[LoadQueue.scala 78:18:@5303.6]
  assign _GEN_200 = 4'he == _T_2022 ? 1'h0 : _GEN_199; // @[LoadQueue.scala 78:18:@5303.6]
  assign _GEN_201 = 4'hf == _T_2022 ? 1'h0 : _GEN_200; // @[LoadQueue.scala 78:18:@5303.6]
  assign _GEN_202 = initBits_5 ? _GEN_185 : offsetQ_5; // @[LoadQueue.scala 76:25:@5289.4]
  assign _GEN_203 = initBits_5 ? _GEN_201 : portQ_5; // @[LoadQueue.scala 76:25:@5289.4]
  assign _T_2040 = _T_1781[3:0]; // @[:@5311.6]
  assign _GEN_205 = 4'h1 == _T_2040 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_206 = 4'h2 == _T_2040 ? io_bbLoadOffsets_2 : _GEN_205; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_207 = 4'h3 == _T_2040 ? io_bbLoadOffsets_3 : _GEN_206; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_208 = 4'h4 == _T_2040 ? io_bbLoadOffsets_4 : _GEN_207; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_209 = 4'h5 == _T_2040 ? io_bbLoadOffsets_5 : _GEN_208; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_210 = 4'h6 == _T_2040 ? io_bbLoadOffsets_6 : _GEN_209; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_211 = 4'h7 == _T_2040 ? io_bbLoadOffsets_7 : _GEN_210; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_212 = 4'h8 == _T_2040 ? io_bbLoadOffsets_8 : _GEN_211; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_213 = 4'h9 == _T_2040 ? io_bbLoadOffsets_9 : _GEN_212; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_214 = 4'ha == _T_2040 ? io_bbLoadOffsets_10 : _GEN_213; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_215 = 4'hb == _T_2040 ? io_bbLoadOffsets_11 : _GEN_214; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_216 = 4'hc == _T_2040 ? io_bbLoadOffsets_12 : _GEN_215; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_217 = 4'hd == _T_2040 ? io_bbLoadOffsets_13 : _GEN_216; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_218 = 4'he == _T_2040 ? io_bbLoadOffsets_14 : _GEN_217; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_219 = 4'hf == _T_2040 ? io_bbLoadOffsets_15 : _GEN_218; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_221 = 4'h1 == _T_2040 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@5319.6]
  assign _GEN_222 = 4'h2 == _T_2040 ? 1'h0 : _GEN_221; // @[LoadQueue.scala 78:18:@5319.6]
  assign _GEN_223 = 4'h3 == _T_2040 ? 1'h0 : _GEN_222; // @[LoadQueue.scala 78:18:@5319.6]
  assign _GEN_224 = 4'h4 == _T_2040 ? 1'h0 : _GEN_223; // @[LoadQueue.scala 78:18:@5319.6]
  assign _GEN_225 = 4'h5 == _T_2040 ? 1'h0 : _GEN_224; // @[LoadQueue.scala 78:18:@5319.6]
  assign _GEN_226 = 4'h6 == _T_2040 ? 1'h0 : _GEN_225; // @[LoadQueue.scala 78:18:@5319.6]
  assign _GEN_227 = 4'h7 == _T_2040 ? 1'h0 : _GEN_226; // @[LoadQueue.scala 78:18:@5319.6]
  assign _GEN_228 = 4'h8 == _T_2040 ? 1'h0 : _GEN_227; // @[LoadQueue.scala 78:18:@5319.6]
  assign _GEN_229 = 4'h9 == _T_2040 ? 1'h0 : _GEN_228; // @[LoadQueue.scala 78:18:@5319.6]
  assign _GEN_230 = 4'ha == _T_2040 ? 1'h0 : _GEN_229; // @[LoadQueue.scala 78:18:@5319.6]
  assign _GEN_231 = 4'hb == _T_2040 ? 1'h0 : _GEN_230; // @[LoadQueue.scala 78:18:@5319.6]
  assign _GEN_232 = 4'hc == _T_2040 ? 1'h0 : _GEN_231; // @[LoadQueue.scala 78:18:@5319.6]
  assign _GEN_233 = 4'hd == _T_2040 ? 1'h0 : _GEN_232; // @[LoadQueue.scala 78:18:@5319.6]
  assign _GEN_234 = 4'he == _T_2040 ? 1'h0 : _GEN_233; // @[LoadQueue.scala 78:18:@5319.6]
  assign _GEN_235 = 4'hf == _T_2040 ? 1'h0 : _GEN_234; // @[LoadQueue.scala 78:18:@5319.6]
  assign _GEN_236 = initBits_6 ? _GEN_219 : offsetQ_6; // @[LoadQueue.scala 76:25:@5305.4]
  assign _GEN_237 = initBits_6 ? _GEN_235 : portQ_6; // @[LoadQueue.scala 76:25:@5305.4]
  assign _T_2058 = _T_1790[3:0]; // @[:@5327.6]
  assign _GEN_239 = 4'h1 == _T_2058 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_240 = 4'h2 == _T_2058 ? io_bbLoadOffsets_2 : _GEN_239; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_241 = 4'h3 == _T_2058 ? io_bbLoadOffsets_3 : _GEN_240; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_242 = 4'h4 == _T_2058 ? io_bbLoadOffsets_4 : _GEN_241; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_243 = 4'h5 == _T_2058 ? io_bbLoadOffsets_5 : _GEN_242; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_244 = 4'h6 == _T_2058 ? io_bbLoadOffsets_6 : _GEN_243; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_245 = 4'h7 == _T_2058 ? io_bbLoadOffsets_7 : _GEN_244; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_246 = 4'h8 == _T_2058 ? io_bbLoadOffsets_8 : _GEN_245; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_247 = 4'h9 == _T_2058 ? io_bbLoadOffsets_9 : _GEN_246; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_248 = 4'ha == _T_2058 ? io_bbLoadOffsets_10 : _GEN_247; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_249 = 4'hb == _T_2058 ? io_bbLoadOffsets_11 : _GEN_248; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_250 = 4'hc == _T_2058 ? io_bbLoadOffsets_12 : _GEN_249; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_251 = 4'hd == _T_2058 ? io_bbLoadOffsets_13 : _GEN_250; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_252 = 4'he == _T_2058 ? io_bbLoadOffsets_14 : _GEN_251; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_253 = 4'hf == _T_2058 ? io_bbLoadOffsets_15 : _GEN_252; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_255 = 4'h1 == _T_2058 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@5335.6]
  assign _GEN_256 = 4'h2 == _T_2058 ? 1'h0 : _GEN_255; // @[LoadQueue.scala 78:18:@5335.6]
  assign _GEN_257 = 4'h3 == _T_2058 ? 1'h0 : _GEN_256; // @[LoadQueue.scala 78:18:@5335.6]
  assign _GEN_258 = 4'h4 == _T_2058 ? 1'h0 : _GEN_257; // @[LoadQueue.scala 78:18:@5335.6]
  assign _GEN_259 = 4'h5 == _T_2058 ? 1'h0 : _GEN_258; // @[LoadQueue.scala 78:18:@5335.6]
  assign _GEN_260 = 4'h6 == _T_2058 ? 1'h0 : _GEN_259; // @[LoadQueue.scala 78:18:@5335.6]
  assign _GEN_261 = 4'h7 == _T_2058 ? 1'h0 : _GEN_260; // @[LoadQueue.scala 78:18:@5335.6]
  assign _GEN_262 = 4'h8 == _T_2058 ? 1'h0 : _GEN_261; // @[LoadQueue.scala 78:18:@5335.6]
  assign _GEN_263 = 4'h9 == _T_2058 ? 1'h0 : _GEN_262; // @[LoadQueue.scala 78:18:@5335.6]
  assign _GEN_264 = 4'ha == _T_2058 ? 1'h0 : _GEN_263; // @[LoadQueue.scala 78:18:@5335.6]
  assign _GEN_265 = 4'hb == _T_2058 ? 1'h0 : _GEN_264; // @[LoadQueue.scala 78:18:@5335.6]
  assign _GEN_266 = 4'hc == _T_2058 ? 1'h0 : _GEN_265; // @[LoadQueue.scala 78:18:@5335.6]
  assign _GEN_267 = 4'hd == _T_2058 ? 1'h0 : _GEN_266; // @[LoadQueue.scala 78:18:@5335.6]
  assign _GEN_268 = 4'he == _T_2058 ? 1'h0 : _GEN_267; // @[LoadQueue.scala 78:18:@5335.6]
  assign _GEN_269 = 4'hf == _T_2058 ? 1'h0 : _GEN_268; // @[LoadQueue.scala 78:18:@5335.6]
  assign _GEN_270 = initBits_7 ? _GEN_253 : offsetQ_7; // @[LoadQueue.scala 76:25:@5321.4]
  assign _GEN_271 = initBits_7 ? _GEN_269 : portQ_7; // @[LoadQueue.scala 76:25:@5321.4]
  assign _T_2076 = _T_1799[3:0]; // @[:@5343.6]
  assign _GEN_273 = 4'h1 == _T_2076 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_274 = 4'h2 == _T_2076 ? io_bbLoadOffsets_2 : _GEN_273; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_275 = 4'h3 == _T_2076 ? io_bbLoadOffsets_3 : _GEN_274; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_276 = 4'h4 == _T_2076 ? io_bbLoadOffsets_4 : _GEN_275; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_277 = 4'h5 == _T_2076 ? io_bbLoadOffsets_5 : _GEN_276; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_278 = 4'h6 == _T_2076 ? io_bbLoadOffsets_6 : _GEN_277; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_279 = 4'h7 == _T_2076 ? io_bbLoadOffsets_7 : _GEN_278; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_280 = 4'h8 == _T_2076 ? io_bbLoadOffsets_8 : _GEN_279; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_281 = 4'h9 == _T_2076 ? io_bbLoadOffsets_9 : _GEN_280; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_282 = 4'ha == _T_2076 ? io_bbLoadOffsets_10 : _GEN_281; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_283 = 4'hb == _T_2076 ? io_bbLoadOffsets_11 : _GEN_282; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_284 = 4'hc == _T_2076 ? io_bbLoadOffsets_12 : _GEN_283; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_285 = 4'hd == _T_2076 ? io_bbLoadOffsets_13 : _GEN_284; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_286 = 4'he == _T_2076 ? io_bbLoadOffsets_14 : _GEN_285; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_287 = 4'hf == _T_2076 ? io_bbLoadOffsets_15 : _GEN_286; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_289 = 4'h1 == _T_2076 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@5351.6]
  assign _GEN_290 = 4'h2 == _T_2076 ? 1'h0 : _GEN_289; // @[LoadQueue.scala 78:18:@5351.6]
  assign _GEN_291 = 4'h3 == _T_2076 ? 1'h0 : _GEN_290; // @[LoadQueue.scala 78:18:@5351.6]
  assign _GEN_292 = 4'h4 == _T_2076 ? 1'h0 : _GEN_291; // @[LoadQueue.scala 78:18:@5351.6]
  assign _GEN_293 = 4'h5 == _T_2076 ? 1'h0 : _GEN_292; // @[LoadQueue.scala 78:18:@5351.6]
  assign _GEN_294 = 4'h6 == _T_2076 ? 1'h0 : _GEN_293; // @[LoadQueue.scala 78:18:@5351.6]
  assign _GEN_295 = 4'h7 == _T_2076 ? 1'h0 : _GEN_294; // @[LoadQueue.scala 78:18:@5351.6]
  assign _GEN_296 = 4'h8 == _T_2076 ? 1'h0 : _GEN_295; // @[LoadQueue.scala 78:18:@5351.6]
  assign _GEN_297 = 4'h9 == _T_2076 ? 1'h0 : _GEN_296; // @[LoadQueue.scala 78:18:@5351.6]
  assign _GEN_298 = 4'ha == _T_2076 ? 1'h0 : _GEN_297; // @[LoadQueue.scala 78:18:@5351.6]
  assign _GEN_299 = 4'hb == _T_2076 ? 1'h0 : _GEN_298; // @[LoadQueue.scala 78:18:@5351.6]
  assign _GEN_300 = 4'hc == _T_2076 ? 1'h0 : _GEN_299; // @[LoadQueue.scala 78:18:@5351.6]
  assign _GEN_301 = 4'hd == _T_2076 ? 1'h0 : _GEN_300; // @[LoadQueue.scala 78:18:@5351.6]
  assign _GEN_302 = 4'he == _T_2076 ? 1'h0 : _GEN_301; // @[LoadQueue.scala 78:18:@5351.6]
  assign _GEN_303 = 4'hf == _T_2076 ? 1'h0 : _GEN_302; // @[LoadQueue.scala 78:18:@5351.6]
  assign _GEN_304 = initBits_8 ? _GEN_287 : offsetQ_8; // @[LoadQueue.scala 76:25:@5337.4]
  assign _GEN_305 = initBits_8 ? _GEN_303 : portQ_8; // @[LoadQueue.scala 76:25:@5337.4]
  assign _T_2094 = _T_1808[3:0]; // @[:@5359.6]
  assign _GEN_307 = 4'h1 == _T_2094 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_308 = 4'h2 == _T_2094 ? io_bbLoadOffsets_2 : _GEN_307; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_309 = 4'h3 == _T_2094 ? io_bbLoadOffsets_3 : _GEN_308; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_310 = 4'h4 == _T_2094 ? io_bbLoadOffsets_4 : _GEN_309; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_311 = 4'h5 == _T_2094 ? io_bbLoadOffsets_5 : _GEN_310; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_312 = 4'h6 == _T_2094 ? io_bbLoadOffsets_6 : _GEN_311; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_313 = 4'h7 == _T_2094 ? io_bbLoadOffsets_7 : _GEN_312; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_314 = 4'h8 == _T_2094 ? io_bbLoadOffsets_8 : _GEN_313; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_315 = 4'h9 == _T_2094 ? io_bbLoadOffsets_9 : _GEN_314; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_316 = 4'ha == _T_2094 ? io_bbLoadOffsets_10 : _GEN_315; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_317 = 4'hb == _T_2094 ? io_bbLoadOffsets_11 : _GEN_316; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_318 = 4'hc == _T_2094 ? io_bbLoadOffsets_12 : _GEN_317; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_319 = 4'hd == _T_2094 ? io_bbLoadOffsets_13 : _GEN_318; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_320 = 4'he == _T_2094 ? io_bbLoadOffsets_14 : _GEN_319; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_321 = 4'hf == _T_2094 ? io_bbLoadOffsets_15 : _GEN_320; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_323 = 4'h1 == _T_2094 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@5367.6]
  assign _GEN_324 = 4'h2 == _T_2094 ? 1'h0 : _GEN_323; // @[LoadQueue.scala 78:18:@5367.6]
  assign _GEN_325 = 4'h3 == _T_2094 ? 1'h0 : _GEN_324; // @[LoadQueue.scala 78:18:@5367.6]
  assign _GEN_326 = 4'h4 == _T_2094 ? 1'h0 : _GEN_325; // @[LoadQueue.scala 78:18:@5367.6]
  assign _GEN_327 = 4'h5 == _T_2094 ? 1'h0 : _GEN_326; // @[LoadQueue.scala 78:18:@5367.6]
  assign _GEN_328 = 4'h6 == _T_2094 ? 1'h0 : _GEN_327; // @[LoadQueue.scala 78:18:@5367.6]
  assign _GEN_329 = 4'h7 == _T_2094 ? 1'h0 : _GEN_328; // @[LoadQueue.scala 78:18:@5367.6]
  assign _GEN_330 = 4'h8 == _T_2094 ? 1'h0 : _GEN_329; // @[LoadQueue.scala 78:18:@5367.6]
  assign _GEN_331 = 4'h9 == _T_2094 ? 1'h0 : _GEN_330; // @[LoadQueue.scala 78:18:@5367.6]
  assign _GEN_332 = 4'ha == _T_2094 ? 1'h0 : _GEN_331; // @[LoadQueue.scala 78:18:@5367.6]
  assign _GEN_333 = 4'hb == _T_2094 ? 1'h0 : _GEN_332; // @[LoadQueue.scala 78:18:@5367.6]
  assign _GEN_334 = 4'hc == _T_2094 ? 1'h0 : _GEN_333; // @[LoadQueue.scala 78:18:@5367.6]
  assign _GEN_335 = 4'hd == _T_2094 ? 1'h0 : _GEN_334; // @[LoadQueue.scala 78:18:@5367.6]
  assign _GEN_336 = 4'he == _T_2094 ? 1'h0 : _GEN_335; // @[LoadQueue.scala 78:18:@5367.6]
  assign _GEN_337 = 4'hf == _T_2094 ? 1'h0 : _GEN_336; // @[LoadQueue.scala 78:18:@5367.6]
  assign _GEN_338 = initBits_9 ? _GEN_321 : offsetQ_9; // @[LoadQueue.scala 76:25:@5353.4]
  assign _GEN_339 = initBits_9 ? _GEN_337 : portQ_9; // @[LoadQueue.scala 76:25:@5353.4]
  assign _T_2112 = _T_1817[3:0]; // @[:@5375.6]
  assign _GEN_341 = 4'h1 == _T_2112 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_342 = 4'h2 == _T_2112 ? io_bbLoadOffsets_2 : _GEN_341; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_343 = 4'h3 == _T_2112 ? io_bbLoadOffsets_3 : _GEN_342; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_344 = 4'h4 == _T_2112 ? io_bbLoadOffsets_4 : _GEN_343; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_345 = 4'h5 == _T_2112 ? io_bbLoadOffsets_5 : _GEN_344; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_346 = 4'h6 == _T_2112 ? io_bbLoadOffsets_6 : _GEN_345; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_347 = 4'h7 == _T_2112 ? io_bbLoadOffsets_7 : _GEN_346; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_348 = 4'h8 == _T_2112 ? io_bbLoadOffsets_8 : _GEN_347; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_349 = 4'h9 == _T_2112 ? io_bbLoadOffsets_9 : _GEN_348; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_350 = 4'ha == _T_2112 ? io_bbLoadOffsets_10 : _GEN_349; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_351 = 4'hb == _T_2112 ? io_bbLoadOffsets_11 : _GEN_350; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_352 = 4'hc == _T_2112 ? io_bbLoadOffsets_12 : _GEN_351; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_353 = 4'hd == _T_2112 ? io_bbLoadOffsets_13 : _GEN_352; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_354 = 4'he == _T_2112 ? io_bbLoadOffsets_14 : _GEN_353; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_355 = 4'hf == _T_2112 ? io_bbLoadOffsets_15 : _GEN_354; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_357 = 4'h1 == _T_2112 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@5383.6]
  assign _GEN_358 = 4'h2 == _T_2112 ? 1'h0 : _GEN_357; // @[LoadQueue.scala 78:18:@5383.6]
  assign _GEN_359 = 4'h3 == _T_2112 ? 1'h0 : _GEN_358; // @[LoadQueue.scala 78:18:@5383.6]
  assign _GEN_360 = 4'h4 == _T_2112 ? 1'h0 : _GEN_359; // @[LoadQueue.scala 78:18:@5383.6]
  assign _GEN_361 = 4'h5 == _T_2112 ? 1'h0 : _GEN_360; // @[LoadQueue.scala 78:18:@5383.6]
  assign _GEN_362 = 4'h6 == _T_2112 ? 1'h0 : _GEN_361; // @[LoadQueue.scala 78:18:@5383.6]
  assign _GEN_363 = 4'h7 == _T_2112 ? 1'h0 : _GEN_362; // @[LoadQueue.scala 78:18:@5383.6]
  assign _GEN_364 = 4'h8 == _T_2112 ? 1'h0 : _GEN_363; // @[LoadQueue.scala 78:18:@5383.6]
  assign _GEN_365 = 4'h9 == _T_2112 ? 1'h0 : _GEN_364; // @[LoadQueue.scala 78:18:@5383.6]
  assign _GEN_366 = 4'ha == _T_2112 ? 1'h0 : _GEN_365; // @[LoadQueue.scala 78:18:@5383.6]
  assign _GEN_367 = 4'hb == _T_2112 ? 1'h0 : _GEN_366; // @[LoadQueue.scala 78:18:@5383.6]
  assign _GEN_368 = 4'hc == _T_2112 ? 1'h0 : _GEN_367; // @[LoadQueue.scala 78:18:@5383.6]
  assign _GEN_369 = 4'hd == _T_2112 ? 1'h0 : _GEN_368; // @[LoadQueue.scala 78:18:@5383.6]
  assign _GEN_370 = 4'he == _T_2112 ? 1'h0 : _GEN_369; // @[LoadQueue.scala 78:18:@5383.6]
  assign _GEN_371 = 4'hf == _T_2112 ? 1'h0 : _GEN_370; // @[LoadQueue.scala 78:18:@5383.6]
  assign _GEN_372 = initBits_10 ? _GEN_355 : offsetQ_10; // @[LoadQueue.scala 76:25:@5369.4]
  assign _GEN_373 = initBits_10 ? _GEN_371 : portQ_10; // @[LoadQueue.scala 76:25:@5369.4]
  assign _T_2130 = _T_1826[3:0]; // @[:@5391.6]
  assign _GEN_375 = 4'h1 == _T_2130 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_376 = 4'h2 == _T_2130 ? io_bbLoadOffsets_2 : _GEN_375; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_377 = 4'h3 == _T_2130 ? io_bbLoadOffsets_3 : _GEN_376; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_378 = 4'h4 == _T_2130 ? io_bbLoadOffsets_4 : _GEN_377; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_379 = 4'h5 == _T_2130 ? io_bbLoadOffsets_5 : _GEN_378; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_380 = 4'h6 == _T_2130 ? io_bbLoadOffsets_6 : _GEN_379; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_381 = 4'h7 == _T_2130 ? io_bbLoadOffsets_7 : _GEN_380; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_382 = 4'h8 == _T_2130 ? io_bbLoadOffsets_8 : _GEN_381; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_383 = 4'h9 == _T_2130 ? io_bbLoadOffsets_9 : _GEN_382; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_384 = 4'ha == _T_2130 ? io_bbLoadOffsets_10 : _GEN_383; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_385 = 4'hb == _T_2130 ? io_bbLoadOffsets_11 : _GEN_384; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_386 = 4'hc == _T_2130 ? io_bbLoadOffsets_12 : _GEN_385; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_387 = 4'hd == _T_2130 ? io_bbLoadOffsets_13 : _GEN_386; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_388 = 4'he == _T_2130 ? io_bbLoadOffsets_14 : _GEN_387; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_389 = 4'hf == _T_2130 ? io_bbLoadOffsets_15 : _GEN_388; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_391 = 4'h1 == _T_2130 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@5399.6]
  assign _GEN_392 = 4'h2 == _T_2130 ? 1'h0 : _GEN_391; // @[LoadQueue.scala 78:18:@5399.6]
  assign _GEN_393 = 4'h3 == _T_2130 ? 1'h0 : _GEN_392; // @[LoadQueue.scala 78:18:@5399.6]
  assign _GEN_394 = 4'h4 == _T_2130 ? 1'h0 : _GEN_393; // @[LoadQueue.scala 78:18:@5399.6]
  assign _GEN_395 = 4'h5 == _T_2130 ? 1'h0 : _GEN_394; // @[LoadQueue.scala 78:18:@5399.6]
  assign _GEN_396 = 4'h6 == _T_2130 ? 1'h0 : _GEN_395; // @[LoadQueue.scala 78:18:@5399.6]
  assign _GEN_397 = 4'h7 == _T_2130 ? 1'h0 : _GEN_396; // @[LoadQueue.scala 78:18:@5399.6]
  assign _GEN_398 = 4'h8 == _T_2130 ? 1'h0 : _GEN_397; // @[LoadQueue.scala 78:18:@5399.6]
  assign _GEN_399 = 4'h9 == _T_2130 ? 1'h0 : _GEN_398; // @[LoadQueue.scala 78:18:@5399.6]
  assign _GEN_400 = 4'ha == _T_2130 ? 1'h0 : _GEN_399; // @[LoadQueue.scala 78:18:@5399.6]
  assign _GEN_401 = 4'hb == _T_2130 ? 1'h0 : _GEN_400; // @[LoadQueue.scala 78:18:@5399.6]
  assign _GEN_402 = 4'hc == _T_2130 ? 1'h0 : _GEN_401; // @[LoadQueue.scala 78:18:@5399.6]
  assign _GEN_403 = 4'hd == _T_2130 ? 1'h0 : _GEN_402; // @[LoadQueue.scala 78:18:@5399.6]
  assign _GEN_404 = 4'he == _T_2130 ? 1'h0 : _GEN_403; // @[LoadQueue.scala 78:18:@5399.6]
  assign _GEN_405 = 4'hf == _T_2130 ? 1'h0 : _GEN_404; // @[LoadQueue.scala 78:18:@5399.6]
  assign _GEN_406 = initBits_11 ? _GEN_389 : offsetQ_11; // @[LoadQueue.scala 76:25:@5385.4]
  assign _GEN_407 = initBits_11 ? _GEN_405 : portQ_11; // @[LoadQueue.scala 76:25:@5385.4]
  assign _T_2148 = _T_1835[3:0]; // @[:@5407.6]
  assign _GEN_409 = 4'h1 == _T_2148 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_410 = 4'h2 == _T_2148 ? io_bbLoadOffsets_2 : _GEN_409; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_411 = 4'h3 == _T_2148 ? io_bbLoadOffsets_3 : _GEN_410; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_412 = 4'h4 == _T_2148 ? io_bbLoadOffsets_4 : _GEN_411; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_413 = 4'h5 == _T_2148 ? io_bbLoadOffsets_5 : _GEN_412; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_414 = 4'h6 == _T_2148 ? io_bbLoadOffsets_6 : _GEN_413; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_415 = 4'h7 == _T_2148 ? io_bbLoadOffsets_7 : _GEN_414; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_416 = 4'h8 == _T_2148 ? io_bbLoadOffsets_8 : _GEN_415; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_417 = 4'h9 == _T_2148 ? io_bbLoadOffsets_9 : _GEN_416; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_418 = 4'ha == _T_2148 ? io_bbLoadOffsets_10 : _GEN_417; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_419 = 4'hb == _T_2148 ? io_bbLoadOffsets_11 : _GEN_418; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_420 = 4'hc == _T_2148 ? io_bbLoadOffsets_12 : _GEN_419; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_421 = 4'hd == _T_2148 ? io_bbLoadOffsets_13 : _GEN_420; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_422 = 4'he == _T_2148 ? io_bbLoadOffsets_14 : _GEN_421; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_423 = 4'hf == _T_2148 ? io_bbLoadOffsets_15 : _GEN_422; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_425 = 4'h1 == _T_2148 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@5415.6]
  assign _GEN_426 = 4'h2 == _T_2148 ? 1'h0 : _GEN_425; // @[LoadQueue.scala 78:18:@5415.6]
  assign _GEN_427 = 4'h3 == _T_2148 ? 1'h0 : _GEN_426; // @[LoadQueue.scala 78:18:@5415.6]
  assign _GEN_428 = 4'h4 == _T_2148 ? 1'h0 : _GEN_427; // @[LoadQueue.scala 78:18:@5415.6]
  assign _GEN_429 = 4'h5 == _T_2148 ? 1'h0 : _GEN_428; // @[LoadQueue.scala 78:18:@5415.6]
  assign _GEN_430 = 4'h6 == _T_2148 ? 1'h0 : _GEN_429; // @[LoadQueue.scala 78:18:@5415.6]
  assign _GEN_431 = 4'h7 == _T_2148 ? 1'h0 : _GEN_430; // @[LoadQueue.scala 78:18:@5415.6]
  assign _GEN_432 = 4'h8 == _T_2148 ? 1'h0 : _GEN_431; // @[LoadQueue.scala 78:18:@5415.6]
  assign _GEN_433 = 4'h9 == _T_2148 ? 1'h0 : _GEN_432; // @[LoadQueue.scala 78:18:@5415.6]
  assign _GEN_434 = 4'ha == _T_2148 ? 1'h0 : _GEN_433; // @[LoadQueue.scala 78:18:@5415.6]
  assign _GEN_435 = 4'hb == _T_2148 ? 1'h0 : _GEN_434; // @[LoadQueue.scala 78:18:@5415.6]
  assign _GEN_436 = 4'hc == _T_2148 ? 1'h0 : _GEN_435; // @[LoadQueue.scala 78:18:@5415.6]
  assign _GEN_437 = 4'hd == _T_2148 ? 1'h0 : _GEN_436; // @[LoadQueue.scala 78:18:@5415.6]
  assign _GEN_438 = 4'he == _T_2148 ? 1'h0 : _GEN_437; // @[LoadQueue.scala 78:18:@5415.6]
  assign _GEN_439 = 4'hf == _T_2148 ? 1'h0 : _GEN_438; // @[LoadQueue.scala 78:18:@5415.6]
  assign _GEN_440 = initBits_12 ? _GEN_423 : offsetQ_12; // @[LoadQueue.scala 76:25:@5401.4]
  assign _GEN_441 = initBits_12 ? _GEN_439 : portQ_12; // @[LoadQueue.scala 76:25:@5401.4]
  assign _T_2166 = _T_1844[3:0]; // @[:@5423.6]
  assign _GEN_443 = 4'h1 == _T_2166 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_444 = 4'h2 == _T_2166 ? io_bbLoadOffsets_2 : _GEN_443; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_445 = 4'h3 == _T_2166 ? io_bbLoadOffsets_3 : _GEN_444; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_446 = 4'h4 == _T_2166 ? io_bbLoadOffsets_4 : _GEN_445; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_447 = 4'h5 == _T_2166 ? io_bbLoadOffsets_5 : _GEN_446; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_448 = 4'h6 == _T_2166 ? io_bbLoadOffsets_6 : _GEN_447; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_449 = 4'h7 == _T_2166 ? io_bbLoadOffsets_7 : _GEN_448; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_450 = 4'h8 == _T_2166 ? io_bbLoadOffsets_8 : _GEN_449; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_451 = 4'h9 == _T_2166 ? io_bbLoadOffsets_9 : _GEN_450; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_452 = 4'ha == _T_2166 ? io_bbLoadOffsets_10 : _GEN_451; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_453 = 4'hb == _T_2166 ? io_bbLoadOffsets_11 : _GEN_452; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_454 = 4'hc == _T_2166 ? io_bbLoadOffsets_12 : _GEN_453; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_455 = 4'hd == _T_2166 ? io_bbLoadOffsets_13 : _GEN_454; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_456 = 4'he == _T_2166 ? io_bbLoadOffsets_14 : _GEN_455; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_457 = 4'hf == _T_2166 ? io_bbLoadOffsets_15 : _GEN_456; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_459 = 4'h1 == _T_2166 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@5431.6]
  assign _GEN_460 = 4'h2 == _T_2166 ? 1'h0 : _GEN_459; // @[LoadQueue.scala 78:18:@5431.6]
  assign _GEN_461 = 4'h3 == _T_2166 ? 1'h0 : _GEN_460; // @[LoadQueue.scala 78:18:@5431.6]
  assign _GEN_462 = 4'h4 == _T_2166 ? 1'h0 : _GEN_461; // @[LoadQueue.scala 78:18:@5431.6]
  assign _GEN_463 = 4'h5 == _T_2166 ? 1'h0 : _GEN_462; // @[LoadQueue.scala 78:18:@5431.6]
  assign _GEN_464 = 4'h6 == _T_2166 ? 1'h0 : _GEN_463; // @[LoadQueue.scala 78:18:@5431.6]
  assign _GEN_465 = 4'h7 == _T_2166 ? 1'h0 : _GEN_464; // @[LoadQueue.scala 78:18:@5431.6]
  assign _GEN_466 = 4'h8 == _T_2166 ? 1'h0 : _GEN_465; // @[LoadQueue.scala 78:18:@5431.6]
  assign _GEN_467 = 4'h9 == _T_2166 ? 1'h0 : _GEN_466; // @[LoadQueue.scala 78:18:@5431.6]
  assign _GEN_468 = 4'ha == _T_2166 ? 1'h0 : _GEN_467; // @[LoadQueue.scala 78:18:@5431.6]
  assign _GEN_469 = 4'hb == _T_2166 ? 1'h0 : _GEN_468; // @[LoadQueue.scala 78:18:@5431.6]
  assign _GEN_470 = 4'hc == _T_2166 ? 1'h0 : _GEN_469; // @[LoadQueue.scala 78:18:@5431.6]
  assign _GEN_471 = 4'hd == _T_2166 ? 1'h0 : _GEN_470; // @[LoadQueue.scala 78:18:@5431.6]
  assign _GEN_472 = 4'he == _T_2166 ? 1'h0 : _GEN_471; // @[LoadQueue.scala 78:18:@5431.6]
  assign _GEN_473 = 4'hf == _T_2166 ? 1'h0 : _GEN_472; // @[LoadQueue.scala 78:18:@5431.6]
  assign _GEN_474 = initBits_13 ? _GEN_457 : offsetQ_13; // @[LoadQueue.scala 76:25:@5417.4]
  assign _GEN_475 = initBits_13 ? _GEN_473 : portQ_13; // @[LoadQueue.scala 76:25:@5417.4]
  assign _T_2184 = _T_1853[3:0]; // @[:@5439.6]
  assign _GEN_477 = 4'h1 == _T_2184 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_478 = 4'h2 == _T_2184 ? io_bbLoadOffsets_2 : _GEN_477; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_479 = 4'h3 == _T_2184 ? io_bbLoadOffsets_3 : _GEN_478; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_480 = 4'h4 == _T_2184 ? io_bbLoadOffsets_4 : _GEN_479; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_481 = 4'h5 == _T_2184 ? io_bbLoadOffsets_5 : _GEN_480; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_482 = 4'h6 == _T_2184 ? io_bbLoadOffsets_6 : _GEN_481; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_483 = 4'h7 == _T_2184 ? io_bbLoadOffsets_7 : _GEN_482; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_484 = 4'h8 == _T_2184 ? io_bbLoadOffsets_8 : _GEN_483; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_485 = 4'h9 == _T_2184 ? io_bbLoadOffsets_9 : _GEN_484; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_486 = 4'ha == _T_2184 ? io_bbLoadOffsets_10 : _GEN_485; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_487 = 4'hb == _T_2184 ? io_bbLoadOffsets_11 : _GEN_486; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_488 = 4'hc == _T_2184 ? io_bbLoadOffsets_12 : _GEN_487; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_489 = 4'hd == _T_2184 ? io_bbLoadOffsets_13 : _GEN_488; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_490 = 4'he == _T_2184 ? io_bbLoadOffsets_14 : _GEN_489; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_491 = 4'hf == _T_2184 ? io_bbLoadOffsets_15 : _GEN_490; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_493 = 4'h1 == _T_2184 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@5447.6]
  assign _GEN_494 = 4'h2 == _T_2184 ? 1'h0 : _GEN_493; // @[LoadQueue.scala 78:18:@5447.6]
  assign _GEN_495 = 4'h3 == _T_2184 ? 1'h0 : _GEN_494; // @[LoadQueue.scala 78:18:@5447.6]
  assign _GEN_496 = 4'h4 == _T_2184 ? 1'h0 : _GEN_495; // @[LoadQueue.scala 78:18:@5447.6]
  assign _GEN_497 = 4'h5 == _T_2184 ? 1'h0 : _GEN_496; // @[LoadQueue.scala 78:18:@5447.6]
  assign _GEN_498 = 4'h6 == _T_2184 ? 1'h0 : _GEN_497; // @[LoadQueue.scala 78:18:@5447.6]
  assign _GEN_499 = 4'h7 == _T_2184 ? 1'h0 : _GEN_498; // @[LoadQueue.scala 78:18:@5447.6]
  assign _GEN_500 = 4'h8 == _T_2184 ? 1'h0 : _GEN_499; // @[LoadQueue.scala 78:18:@5447.6]
  assign _GEN_501 = 4'h9 == _T_2184 ? 1'h0 : _GEN_500; // @[LoadQueue.scala 78:18:@5447.6]
  assign _GEN_502 = 4'ha == _T_2184 ? 1'h0 : _GEN_501; // @[LoadQueue.scala 78:18:@5447.6]
  assign _GEN_503 = 4'hb == _T_2184 ? 1'h0 : _GEN_502; // @[LoadQueue.scala 78:18:@5447.6]
  assign _GEN_504 = 4'hc == _T_2184 ? 1'h0 : _GEN_503; // @[LoadQueue.scala 78:18:@5447.6]
  assign _GEN_505 = 4'hd == _T_2184 ? 1'h0 : _GEN_504; // @[LoadQueue.scala 78:18:@5447.6]
  assign _GEN_506 = 4'he == _T_2184 ? 1'h0 : _GEN_505; // @[LoadQueue.scala 78:18:@5447.6]
  assign _GEN_507 = 4'hf == _T_2184 ? 1'h0 : _GEN_506; // @[LoadQueue.scala 78:18:@5447.6]
  assign _GEN_508 = initBits_14 ? _GEN_491 : offsetQ_14; // @[LoadQueue.scala 76:25:@5433.4]
  assign _GEN_509 = initBits_14 ? _GEN_507 : portQ_14; // @[LoadQueue.scala 76:25:@5433.4]
  assign _T_2202 = _T_1862[3:0]; // @[:@5455.6]
  assign _GEN_511 = 4'h1 == _T_2202 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_512 = 4'h2 == _T_2202 ? io_bbLoadOffsets_2 : _GEN_511; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_513 = 4'h3 == _T_2202 ? io_bbLoadOffsets_3 : _GEN_512; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_514 = 4'h4 == _T_2202 ? io_bbLoadOffsets_4 : _GEN_513; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_515 = 4'h5 == _T_2202 ? io_bbLoadOffsets_5 : _GEN_514; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_516 = 4'h6 == _T_2202 ? io_bbLoadOffsets_6 : _GEN_515; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_517 = 4'h7 == _T_2202 ? io_bbLoadOffsets_7 : _GEN_516; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_518 = 4'h8 == _T_2202 ? io_bbLoadOffsets_8 : _GEN_517; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_519 = 4'h9 == _T_2202 ? io_bbLoadOffsets_9 : _GEN_518; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_520 = 4'ha == _T_2202 ? io_bbLoadOffsets_10 : _GEN_519; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_521 = 4'hb == _T_2202 ? io_bbLoadOffsets_11 : _GEN_520; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_522 = 4'hc == _T_2202 ? io_bbLoadOffsets_12 : _GEN_521; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_523 = 4'hd == _T_2202 ? io_bbLoadOffsets_13 : _GEN_522; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_524 = 4'he == _T_2202 ? io_bbLoadOffsets_14 : _GEN_523; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_525 = 4'hf == _T_2202 ? io_bbLoadOffsets_15 : _GEN_524; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_527 = 4'h1 == _T_2202 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@5463.6]
  assign _GEN_528 = 4'h2 == _T_2202 ? 1'h0 : _GEN_527; // @[LoadQueue.scala 78:18:@5463.6]
  assign _GEN_529 = 4'h3 == _T_2202 ? 1'h0 : _GEN_528; // @[LoadQueue.scala 78:18:@5463.6]
  assign _GEN_530 = 4'h4 == _T_2202 ? 1'h0 : _GEN_529; // @[LoadQueue.scala 78:18:@5463.6]
  assign _GEN_531 = 4'h5 == _T_2202 ? 1'h0 : _GEN_530; // @[LoadQueue.scala 78:18:@5463.6]
  assign _GEN_532 = 4'h6 == _T_2202 ? 1'h0 : _GEN_531; // @[LoadQueue.scala 78:18:@5463.6]
  assign _GEN_533 = 4'h7 == _T_2202 ? 1'h0 : _GEN_532; // @[LoadQueue.scala 78:18:@5463.6]
  assign _GEN_534 = 4'h8 == _T_2202 ? 1'h0 : _GEN_533; // @[LoadQueue.scala 78:18:@5463.6]
  assign _GEN_535 = 4'h9 == _T_2202 ? 1'h0 : _GEN_534; // @[LoadQueue.scala 78:18:@5463.6]
  assign _GEN_536 = 4'ha == _T_2202 ? 1'h0 : _GEN_535; // @[LoadQueue.scala 78:18:@5463.6]
  assign _GEN_537 = 4'hb == _T_2202 ? 1'h0 : _GEN_536; // @[LoadQueue.scala 78:18:@5463.6]
  assign _GEN_538 = 4'hc == _T_2202 ? 1'h0 : _GEN_537; // @[LoadQueue.scala 78:18:@5463.6]
  assign _GEN_539 = 4'hd == _T_2202 ? 1'h0 : _GEN_538; // @[LoadQueue.scala 78:18:@5463.6]
  assign _GEN_540 = 4'he == _T_2202 ? 1'h0 : _GEN_539; // @[LoadQueue.scala 78:18:@5463.6]
  assign _GEN_541 = 4'hf == _T_2202 ? 1'h0 : _GEN_540; // @[LoadQueue.scala 78:18:@5463.6]
  assign _GEN_542 = initBits_15 ? _GEN_525 : offsetQ_15; // @[LoadQueue.scala 76:25:@5449.4]
  assign _GEN_543 = initBits_15 ? _GEN_541 : portQ_15; // @[LoadQueue.scala 76:25:@5449.4]
  assign _T_2224 = _GEN_15 + 4'h1; // @[util.scala 10:8:@5474.6]
  assign _GEN_272 = _T_2224 % 5'h10; // @[util.scala 10:14:@5475.6]
  assign _T_2225 = _GEN_272[4:0]; // @[util.scala 10:14:@5475.6]
  assign _GEN_2377 = {{1'd0}, io_storeTail}; // @[LoadQueue.scala 97:56:@5476.6]
  assign _T_2226 = _T_2225 == _GEN_2377; // @[LoadQueue.scala 97:56:@5476.6]
  assign _T_2227 = io_storeEmpty & _T_2226; // @[LoadQueue.scala 96:50:@5477.6]
  assign _T_2229 = _T_2227 == 1'h0; // @[LoadQueue.scala 96:34:@5478.6]
  assign _T_2231 = previousStoreHead <= offsetQ_0; // @[LoadQueue.scala 101:36:@5486.8]
  assign _T_2232 = offsetQ_0 < io_storeHead; // @[LoadQueue.scala 101:86:@5487.8]
  assign _T_2233 = _T_2231 & _T_2232; // @[LoadQueue.scala 101:61:@5488.8]
  assign _T_2235 = previousStoreHead > io_storeHead; // @[LoadQueue.scala 103:36:@5493.10]
  assign _T_2236 = io_storeHead <= offsetQ_0; // @[LoadQueue.scala 103:69:@5494.10]
  assign _T_2237 = offsetQ_0 < previousStoreHead; // @[LoadQueue.scala 104:31:@5495.10]
  assign _T_2238 = _T_2236 & _T_2237; // @[LoadQueue.scala 103:94:@5496.10]
  assign _T_2240 = _T_2238 == 1'h0; // @[LoadQueue.scala 103:54:@5497.10]
  assign _T_2241 = _T_2235 & _T_2240; // @[LoadQueue.scala 103:51:@5498.10]
  assign _GEN_560 = _T_2241 ? 1'h0 : checkBits_0; // @[LoadQueue.scala 104:53:@5499.10]
  assign _GEN_561 = _T_2233 ? 1'h0 : _GEN_560; // @[LoadQueue.scala 101:102:@5489.8]
  assign _GEN_562 = io_storeEmpty ? 1'h0 : _GEN_561; // @[LoadQueue.scala 99:27:@5482.6]
  assign _GEN_563 = initBits_0 ? _T_2229 : _GEN_562; // @[LoadQueue.scala 95:34:@5467.4]
  assign _T_2254 = _GEN_49 + 4'h1; // @[util.scala 10:8:@5510.6]
  assign _GEN_288 = _T_2254 % 5'h10; // @[util.scala 10:14:@5511.6]
  assign _T_2255 = _GEN_288[4:0]; // @[util.scala 10:14:@5511.6]
  assign _T_2256 = _T_2255 == _GEN_2377; // @[LoadQueue.scala 97:56:@5512.6]
  assign _T_2257 = io_storeEmpty & _T_2256; // @[LoadQueue.scala 96:50:@5513.6]
  assign _T_2259 = _T_2257 == 1'h0; // @[LoadQueue.scala 96:34:@5514.6]
  assign _T_2261 = previousStoreHead <= offsetQ_1; // @[LoadQueue.scala 101:36:@5522.8]
  assign _T_2262 = offsetQ_1 < io_storeHead; // @[LoadQueue.scala 101:86:@5523.8]
  assign _T_2263 = _T_2261 & _T_2262; // @[LoadQueue.scala 101:61:@5524.8]
  assign _T_2266 = io_storeHead <= offsetQ_1; // @[LoadQueue.scala 103:69:@5530.10]
  assign _T_2267 = offsetQ_1 < previousStoreHead; // @[LoadQueue.scala 104:31:@5531.10]
  assign _T_2268 = _T_2266 & _T_2267; // @[LoadQueue.scala 103:94:@5532.10]
  assign _T_2270 = _T_2268 == 1'h0; // @[LoadQueue.scala 103:54:@5533.10]
  assign _T_2271 = _T_2235 & _T_2270; // @[LoadQueue.scala 103:51:@5534.10]
  assign _GEN_580 = _T_2271 ? 1'h0 : checkBits_1; // @[LoadQueue.scala 104:53:@5535.10]
  assign _GEN_581 = _T_2263 ? 1'h0 : _GEN_580; // @[LoadQueue.scala 101:102:@5525.8]
  assign _GEN_582 = io_storeEmpty ? 1'h0 : _GEN_581; // @[LoadQueue.scala 99:27:@5518.6]
  assign _GEN_583 = initBits_1 ? _T_2259 : _GEN_582; // @[LoadQueue.scala 95:34:@5503.4]
  assign _T_2284 = _GEN_83 + 4'h1; // @[util.scala 10:8:@5546.6]
  assign _GEN_306 = _T_2284 % 5'h10; // @[util.scala 10:14:@5547.6]
  assign _T_2285 = _GEN_306[4:0]; // @[util.scala 10:14:@5547.6]
  assign _T_2286 = _T_2285 == _GEN_2377; // @[LoadQueue.scala 97:56:@5548.6]
  assign _T_2287 = io_storeEmpty & _T_2286; // @[LoadQueue.scala 96:50:@5549.6]
  assign _T_2289 = _T_2287 == 1'h0; // @[LoadQueue.scala 96:34:@5550.6]
  assign _T_2291 = previousStoreHead <= offsetQ_2; // @[LoadQueue.scala 101:36:@5558.8]
  assign _T_2292 = offsetQ_2 < io_storeHead; // @[LoadQueue.scala 101:86:@5559.8]
  assign _T_2293 = _T_2291 & _T_2292; // @[LoadQueue.scala 101:61:@5560.8]
  assign _T_2296 = io_storeHead <= offsetQ_2; // @[LoadQueue.scala 103:69:@5566.10]
  assign _T_2297 = offsetQ_2 < previousStoreHead; // @[LoadQueue.scala 104:31:@5567.10]
  assign _T_2298 = _T_2296 & _T_2297; // @[LoadQueue.scala 103:94:@5568.10]
  assign _T_2300 = _T_2298 == 1'h0; // @[LoadQueue.scala 103:54:@5569.10]
  assign _T_2301 = _T_2235 & _T_2300; // @[LoadQueue.scala 103:51:@5570.10]
  assign _GEN_600 = _T_2301 ? 1'h0 : checkBits_2; // @[LoadQueue.scala 104:53:@5571.10]
  assign _GEN_601 = _T_2293 ? 1'h0 : _GEN_600; // @[LoadQueue.scala 101:102:@5561.8]
  assign _GEN_602 = io_storeEmpty ? 1'h0 : _GEN_601; // @[LoadQueue.scala 99:27:@5554.6]
  assign _GEN_603 = initBits_2 ? _T_2289 : _GEN_602; // @[LoadQueue.scala 95:34:@5539.4]
  assign _T_2314 = _GEN_117 + 4'h1; // @[util.scala 10:8:@5582.6]
  assign _GEN_322 = _T_2314 % 5'h10; // @[util.scala 10:14:@5583.6]
  assign _T_2315 = _GEN_322[4:0]; // @[util.scala 10:14:@5583.6]
  assign _T_2316 = _T_2315 == _GEN_2377; // @[LoadQueue.scala 97:56:@5584.6]
  assign _T_2317 = io_storeEmpty & _T_2316; // @[LoadQueue.scala 96:50:@5585.6]
  assign _T_2319 = _T_2317 == 1'h0; // @[LoadQueue.scala 96:34:@5586.6]
  assign _T_2321 = previousStoreHead <= offsetQ_3; // @[LoadQueue.scala 101:36:@5594.8]
  assign _T_2322 = offsetQ_3 < io_storeHead; // @[LoadQueue.scala 101:86:@5595.8]
  assign _T_2323 = _T_2321 & _T_2322; // @[LoadQueue.scala 101:61:@5596.8]
  assign _T_2326 = io_storeHead <= offsetQ_3; // @[LoadQueue.scala 103:69:@5602.10]
  assign _T_2327 = offsetQ_3 < previousStoreHead; // @[LoadQueue.scala 104:31:@5603.10]
  assign _T_2328 = _T_2326 & _T_2327; // @[LoadQueue.scala 103:94:@5604.10]
  assign _T_2330 = _T_2328 == 1'h0; // @[LoadQueue.scala 103:54:@5605.10]
  assign _T_2331 = _T_2235 & _T_2330; // @[LoadQueue.scala 103:51:@5606.10]
  assign _GEN_620 = _T_2331 ? 1'h0 : checkBits_3; // @[LoadQueue.scala 104:53:@5607.10]
  assign _GEN_621 = _T_2323 ? 1'h0 : _GEN_620; // @[LoadQueue.scala 101:102:@5597.8]
  assign _GEN_622 = io_storeEmpty ? 1'h0 : _GEN_621; // @[LoadQueue.scala 99:27:@5590.6]
  assign _GEN_623 = initBits_3 ? _T_2319 : _GEN_622; // @[LoadQueue.scala 95:34:@5575.4]
  assign _T_2344 = _GEN_151 + 4'h1; // @[util.scala 10:8:@5618.6]
  assign _GEN_340 = _T_2344 % 5'h10; // @[util.scala 10:14:@5619.6]
  assign _T_2345 = _GEN_340[4:0]; // @[util.scala 10:14:@5619.6]
  assign _T_2346 = _T_2345 == _GEN_2377; // @[LoadQueue.scala 97:56:@5620.6]
  assign _T_2347 = io_storeEmpty & _T_2346; // @[LoadQueue.scala 96:50:@5621.6]
  assign _T_2349 = _T_2347 == 1'h0; // @[LoadQueue.scala 96:34:@5622.6]
  assign _T_2351 = previousStoreHead <= offsetQ_4; // @[LoadQueue.scala 101:36:@5630.8]
  assign _T_2352 = offsetQ_4 < io_storeHead; // @[LoadQueue.scala 101:86:@5631.8]
  assign _T_2353 = _T_2351 & _T_2352; // @[LoadQueue.scala 101:61:@5632.8]
  assign _T_2356 = io_storeHead <= offsetQ_4; // @[LoadQueue.scala 103:69:@5638.10]
  assign _T_2357 = offsetQ_4 < previousStoreHead; // @[LoadQueue.scala 104:31:@5639.10]
  assign _T_2358 = _T_2356 & _T_2357; // @[LoadQueue.scala 103:94:@5640.10]
  assign _T_2360 = _T_2358 == 1'h0; // @[LoadQueue.scala 103:54:@5641.10]
  assign _T_2361 = _T_2235 & _T_2360; // @[LoadQueue.scala 103:51:@5642.10]
  assign _GEN_640 = _T_2361 ? 1'h0 : checkBits_4; // @[LoadQueue.scala 104:53:@5643.10]
  assign _GEN_641 = _T_2353 ? 1'h0 : _GEN_640; // @[LoadQueue.scala 101:102:@5633.8]
  assign _GEN_642 = io_storeEmpty ? 1'h0 : _GEN_641; // @[LoadQueue.scala 99:27:@5626.6]
  assign _GEN_643 = initBits_4 ? _T_2349 : _GEN_642; // @[LoadQueue.scala 95:34:@5611.4]
  assign _T_2374 = _GEN_185 + 4'h1; // @[util.scala 10:8:@5654.6]
  assign _GEN_356 = _T_2374 % 5'h10; // @[util.scala 10:14:@5655.6]
  assign _T_2375 = _GEN_356[4:0]; // @[util.scala 10:14:@5655.6]
  assign _T_2376 = _T_2375 == _GEN_2377; // @[LoadQueue.scala 97:56:@5656.6]
  assign _T_2377 = io_storeEmpty & _T_2376; // @[LoadQueue.scala 96:50:@5657.6]
  assign _T_2379 = _T_2377 == 1'h0; // @[LoadQueue.scala 96:34:@5658.6]
  assign _T_2381 = previousStoreHead <= offsetQ_5; // @[LoadQueue.scala 101:36:@5666.8]
  assign _T_2382 = offsetQ_5 < io_storeHead; // @[LoadQueue.scala 101:86:@5667.8]
  assign _T_2383 = _T_2381 & _T_2382; // @[LoadQueue.scala 101:61:@5668.8]
  assign _T_2386 = io_storeHead <= offsetQ_5; // @[LoadQueue.scala 103:69:@5674.10]
  assign _T_2387 = offsetQ_5 < previousStoreHead; // @[LoadQueue.scala 104:31:@5675.10]
  assign _T_2388 = _T_2386 & _T_2387; // @[LoadQueue.scala 103:94:@5676.10]
  assign _T_2390 = _T_2388 == 1'h0; // @[LoadQueue.scala 103:54:@5677.10]
  assign _T_2391 = _T_2235 & _T_2390; // @[LoadQueue.scala 103:51:@5678.10]
  assign _GEN_660 = _T_2391 ? 1'h0 : checkBits_5; // @[LoadQueue.scala 104:53:@5679.10]
  assign _GEN_661 = _T_2383 ? 1'h0 : _GEN_660; // @[LoadQueue.scala 101:102:@5669.8]
  assign _GEN_662 = io_storeEmpty ? 1'h0 : _GEN_661; // @[LoadQueue.scala 99:27:@5662.6]
  assign _GEN_663 = initBits_5 ? _T_2379 : _GEN_662; // @[LoadQueue.scala 95:34:@5647.4]
  assign _T_2404 = _GEN_219 + 4'h1; // @[util.scala 10:8:@5690.6]
  assign _GEN_374 = _T_2404 % 5'h10; // @[util.scala 10:14:@5691.6]
  assign _T_2405 = _GEN_374[4:0]; // @[util.scala 10:14:@5691.6]
  assign _T_2406 = _T_2405 == _GEN_2377; // @[LoadQueue.scala 97:56:@5692.6]
  assign _T_2407 = io_storeEmpty & _T_2406; // @[LoadQueue.scala 96:50:@5693.6]
  assign _T_2409 = _T_2407 == 1'h0; // @[LoadQueue.scala 96:34:@5694.6]
  assign _T_2411 = previousStoreHead <= offsetQ_6; // @[LoadQueue.scala 101:36:@5702.8]
  assign _T_2412 = offsetQ_6 < io_storeHead; // @[LoadQueue.scala 101:86:@5703.8]
  assign _T_2413 = _T_2411 & _T_2412; // @[LoadQueue.scala 101:61:@5704.8]
  assign _T_2416 = io_storeHead <= offsetQ_6; // @[LoadQueue.scala 103:69:@5710.10]
  assign _T_2417 = offsetQ_6 < previousStoreHead; // @[LoadQueue.scala 104:31:@5711.10]
  assign _T_2418 = _T_2416 & _T_2417; // @[LoadQueue.scala 103:94:@5712.10]
  assign _T_2420 = _T_2418 == 1'h0; // @[LoadQueue.scala 103:54:@5713.10]
  assign _T_2421 = _T_2235 & _T_2420; // @[LoadQueue.scala 103:51:@5714.10]
  assign _GEN_680 = _T_2421 ? 1'h0 : checkBits_6; // @[LoadQueue.scala 104:53:@5715.10]
  assign _GEN_681 = _T_2413 ? 1'h0 : _GEN_680; // @[LoadQueue.scala 101:102:@5705.8]
  assign _GEN_682 = io_storeEmpty ? 1'h0 : _GEN_681; // @[LoadQueue.scala 99:27:@5698.6]
  assign _GEN_683 = initBits_6 ? _T_2409 : _GEN_682; // @[LoadQueue.scala 95:34:@5683.4]
  assign _T_2434 = _GEN_253 + 4'h1; // @[util.scala 10:8:@5726.6]
  assign _GEN_390 = _T_2434 % 5'h10; // @[util.scala 10:14:@5727.6]
  assign _T_2435 = _GEN_390[4:0]; // @[util.scala 10:14:@5727.6]
  assign _T_2436 = _T_2435 == _GEN_2377; // @[LoadQueue.scala 97:56:@5728.6]
  assign _T_2437 = io_storeEmpty & _T_2436; // @[LoadQueue.scala 96:50:@5729.6]
  assign _T_2439 = _T_2437 == 1'h0; // @[LoadQueue.scala 96:34:@5730.6]
  assign _T_2441 = previousStoreHead <= offsetQ_7; // @[LoadQueue.scala 101:36:@5738.8]
  assign _T_2442 = offsetQ_7 < io_storeHead; // @[LoadQueue.scala 101:86:@5739.8]
  assign _T_2443 = _T_2441 & _T_2442; // @[LoadQueue.scala 101:61:@5740.8]
  assign _T_2446 = io_storeHead <= offsetQ_7; // @[LoadQueue.scala 103:69:@5746.10]
  assign _T_2447 = offsetQ_7 < previousStoreHead; // @[LoadQueue.scala 104:31:@5747.10]
  assign _T_2448 = _T_2446 & _T_2447; // @[LoadQueue.scala 103:94:@5748.10]
  assign _T_2450 = _T_2448 == 1'h0; // @[LoadQueue.scala 103:54:@5749.10]
  assign _T_2451 = _T_2235 & _T_2450; // @[LoadQueue.scala 103:51:@5750.10]
  assign _GEN_700 = _T_2451 ? 1'h0 : checkBits_7; // @[LoadQueue.scala 104:53:@5751.10]
  assign _GEN_701 = _T_2443 ? 1'h0 : _GEN_700; // @[LoadQueue.scala 101:102:@5741.8]
  assign _GEN_702 = io_storeEmpty ? 1'h0 : _GEN_701; // @[LoadQueue.scala 99:27:@5734.6]
  assign _GEN_703 = initBits_7 ? _T_2439 : _GEN_702; // @[LoadQueue.scala 95:34:@5719.4]
  assign _T_2464 = _GEN_287 + 4'h1; // @[util.scala 10:8:@5762.6]
  assign _GEN_408 = _T_2464 % 5'h10; // @[util.scala 10:14:@5763.6]
  assign _T_2465 = _GEN_408[4:0]; // @[util.scala 10:14:@5763.6]
  assign _T_2466 = _T_2465 == _GEN_2377; // @[LoadQueue.scala 97:56:@5764.6]
  assign _T_2467 = io_storeEmpty & _T_2466; // @[LoadQueue.scala 96:50:@5765.6]
  assign _T_2469 = _T_2467 == 1'h0; // @[LoadQueue.scala 96:34:@5766.6]
  assign _T_2471 = previousStoreHead <= offsetQ_8; // @[LoadQueue.scala 101:36:@5774.8]
  assign _T_2472 = offsetQ_8 < io_storeHead; // @[LoadQueue.scala 101:86:@5775.8]
  assign _T_2473 = _T_2471 & _T_2472; // @[LoadQueue.scala 101:61:@5776.8]
  assign _T_2476 = io_storeHead <= offsetQ_8; // @[LoadQueue.scala 103:69:@5782.10]
  assign _T_2477 = offsetQ_8 < previousStoreHead; // @[LoadQueue.scala 104:31:@5783.10]
  assign _T_2478 = _T_2476 & _T_2477; // @[LoadQueue.scala 103:94:@5784.10]
  assign _T_2480 = _T_2478 == 1'h0; // @[LoadQueue.scala 103:54:@5785.10]
  assign _T_2481 = _T_2235 & _T_2480; // @[LoadQueue.scala 103:51:@5786.10]
  assign _GEN_720 = _T_2481 ? 1'h0 : checkBits_8; // @[LoadQueue.scala 104:53:@5787.10]
  assign _GEN_721 = _T_2473 ? 1'h0 : _GEN_720; // @[LoadQueue.scala 101:102:@5777.8]
  assign _GEN_722 = io_storeEmpty ? 1'h0 : _GEN_721; // @[LoadQueue.scala 99:27:@5770.6]
  assign _GEN_723 = initBits_8 ? _T_2469 : _GEN_722; // @[LoadQueue.scala 95:34:@5755.4]
  assign _T_2494 = _GEN_321 + 4'h1; // @[util.scala 10:8:@5798.6]
  assign _GEN_424 = _T_2494 % 5'h10; // @[util.scala 10:14:@5799.6]
  assign _T_2495 = _GEN_424[4:0]; // @[util.scala 10:14:@5799.6]
  assign _T_2496 = _T_2495 == _GEN_2377; // @[LoadQueue.scala 97:56:@5800.6]
  assign _T_2497 = io_storeEmpty & _T_2496; // @[LoadQueue.scala 96:50:@5801.6]
  assign _T_2499 = _T_2497 == 1'h0; // @[LoadQueue.scala 96:34:@5802.6]
  assign _T_2501 = previousStoreHead <= offsetQ_9; // @[LoadQueue.scala 101:36:@5810.8]
  assign _T_2502 = offsetQ_9 < io_storeHead; // @[LoadQueue.scala 101:86:@5811.8]
  assign _T_2503 = _T_2501 & _T_2502; // @[LoadQueue.scala 101:61:@5812.8]
  assign _T_2506 = io_storeHead <= offsetQ_9; // @[LoadQueue.scala 103:69:@5818.10]
  assign _T_2507 = offsetQ_9 < previousStoreHead; // @[LoadQueue.scala 104:31:@5819.10]
  assign _T_2508 = _T_2506 & _T_2507; // @[LoadQueue.scala 103:94:@5820.10]
  assign _T_2510 = _T_2508 == 1'h0; // @[LoadQueue.scala 103:54:@5821.10]
  assign _T_2511 = _T_2235 & _T_2510; // @[LoadQueue.scala 103:51:@5822.10]
  assign _GEN_740 = _T_2511 ? 1'h0 : checkBits_9; // @[LoadQueue.scala 104:53:@5823.10]
  assign _GEN_741 = _T_2503 ? 1'h0 : _GEN_740; // @[LoadQueue.scala 101:102:@5813.8]
  assign _GEN_742 = io_storeEmpty ? 1'h0 : _GEN_741; // @[LoadQueue.scala 99:27:@5806.6]
  assign _GEN_743 = initBits_9 ? _T_2499 : _GEN_742; // @[LoadQueue.scala 95:34:@5791.4]
  assign _T_2524 = _GEN_355 + 4'h1; // @[util.scala 10:8:@5834.6]
  assign _GEN_442 = _T_2524 % 5'h10; // @[util.scala 10:14:@5835.6]
  assign _T_2525 = _GEN_442[4:0]; // @[util.scala 10:14:@5835.6]
  assign _T_2526 = _T_2525 == _GEN_2377; // @[LoadQueue.scala 97:56:@5836.6]
  assign _T_2527 = io_storeEmpty & _T_2526; // @[LoadQueue.scala 96:50:@5837.6]
  assign _T_2529 = _T_2527 == 1'h0; // @[LoadQueue.scala 96:34:@5838.6]
  assign _T_2531 = previousStoreHead <= offsetQ_10; // @[LoadQueue.scala 101:36:@5846.8]
  assign _T_2532 = offsetQ_10 < io_storeHead; // @[LoadQueue.scala 101:86:@5847.8]
  assign _T_2533 = _T_2531 & _T_2532; // @[LoadQueue.scala 101:61:@5848.8]
  assign _T_2536 = io_storeHead <= offsetQ_10; // @[LoadQueue.scala 103:69:@5854.10]
  assign _T_2537 = offsetQ_10 < previousStoreHead; // @[LoadQueue.scala 104:31:@5855.10]
  assign _T_2538 = _T_2536 & _T_2537; // @[LoadQueue.scala 103:94:@5856.10]
  assign _T_2540 = _T_2538 == 1'h0; // @[LoadQueue.scala 103:54:@5857.10]
  assign _T_2541 = _T_2235 & _T_2540; // @[LoadQueue.scala 103:51:@5858.10]
  assign _GEN_760 = _T_2541 ? 1'h0 : checkBits_10; // @[LoadQueue.scala 104:53:@5859.10]
  assign _GEN_761 = _T_2533 ? 1'h0 : _GEN_760; // @[LoadQueue.scala 101:102:@5849.8]
  assign _GEN_762 = io_storeEmpty ? 1'h0 : _GEN_761; // @[LoadQueue.scala 99:27:@5842.6]
  assign _GEN_763 = initBits_10 ? _T_2529 : _GEN_762; // @[LoadQueue.scala 95:34:@5827.4]
  assign _T_2554 = _GEN_389 + 4'h1; // @[util.scala 10:8:@5870.6]
  assign _GEN_458 = _T_2554 % 5'h10; // @[util.scala 10:14:@5871.6]
  assign _T_2555 = _GEN_458[4:0]; // @[util.scala 10:14:@5871.6]
  assign _T_2556 = _T_2555 == _GEN_2377; // @[LoadQueue.scala 97:56:@5872.6]
  assign _T_2557 = io_storeEmpty & _T_2556; // @[LoadQueue.scala 96:50:@5873.6]
  assign _T_2559 = _T_2557 == 1'h0; // @[LoadQueue.scala 96:34:@5874.6]
  assign _T_2561 = previousStoreHead <= offsetQ_11; // @[LoadQueue.scala 101:36:@5882.8]
  assign _T_2562 = offsetQ_11 < io_storeHead; // @[LoadQueue.scala 101:86:@5883.8]
  assign _T_2563 = _T_2561 & _T_2562; // @[LoadQueue.scala 101:61:@5884.8]
  assign _T_2566 = io_storeHead <= offsetQ_11; // @[LoadQueue.scala 103:69:@5890.10]
  assign _T_2567 = offsetQ_11 < previousStoreHead; // @[LoadQueue.scala 104:31:@5891.10]
  assign _T_2568 = _T_2566 & _T_2567; // @[LoadQueue.scala 103:94:@5892.10]
  assign _T_2570 = _T_2568 == 1'h0; // @[LoadQueue.scala 103:54:@5893.10]
  assign _T_2571 = _T_2235 & _T_2570; // @[LoadQueue.scala 103:51:@5894.10]
  assign _GEN_780 = _T_2571 ? 1'h0 : checkBits_11; // @[LoadQueue.scala 104:53:@5895.10]
  assign _GEN_781 = _T_2563 ? 1'h0 : _GEN_780; // @[LoadQueue.scala 101:102:@5885.8]
  assign _GEN_782 = io_storeEmpty ? 1'h0 : _GEN_781; // @[LoadQueue.scala 99:27:@5878.6]
  assign _GEN_783 = initBits_11 ? _T_2559 : _GEN_782; // @[LoadQueue.scala 95:34:@5863.4]
  assign _T_2584 = _GEN_423 + 4'h1; // @[util.scala 10:8:@5906.6]
  assign _GEN_476 = _T_2584 % 5'h10; // @[util.scala 10:14:@5907.6]
  assign _T_2585 = _GEN_476[4:0]; // @[util.scala 10:14:@5907.6]
  assign _T_2586 = _T_2585 == _GEN_2377; // @[LoadQueue.scala 97:56:@5908.6]
  assign _T_2587 = io_storeEmpty & _T_2586; // @[LoadQueue.scala 96:50:@5909.6]
  assign _T_2589 = _T_2587 == 1'h0; // @[LoadQueue.scala 96:34:@5910.6]
  assign _T_2591 = previousStoreHead <= offsetQ_12; // @[LoadQueue.scala 101:36:@5918.8]
  assign _T_2592 = offsetQ_12 < io_storeHead; // @[LoadQueue.scala 101:86:@5919.8]
  assign _T_2593 = _T_2591 & _T_2592; // @[LoadQueue.scala 101:61:@5920.8]
  assign _T_2596 = io_storeHead <= offsetQ_12; // @[LoadQueue.scala 103:69:@5926.10]
  assign _T_2597 = offsetQ_12 < previousStoreHead; // @[LoadQueue.scala 104:31:@5927.10]
  assign _T_2598 = _T_2596 & _T_2597; // @[LoadQueue.scala 103:94:@5928.10]
  assign _T_2600 = _T_2598 == 1'h0; // @[LoadQueue.scala 103:54:@5929.10]
  assign _T_2601 = _T_2235 & _T_2600; // @[LoadQueue.scala 103:51:@5930.10]
  assign _GEN_800 = _T_2601 ? 1'h0 : checkBits_12; // @[LoadQueue.scala 104:53:@5931.10]
  assign _GEN_801 = _T_2593 ? 1'h0 : _GEN_800; // @[LoadQueue.scala 101:102:@5921.8]
  assign _GEN_802 = io_storeEmpty ? 1'h0 : _GEN_801; // @[LoadQueue.scala 99:27:@5914.6]
  assign _GEN_803 = initBits_12 ? _T_2589 : _GEN_802; // @[LoadQueue.scala 95:34:@5899.4]
  assign _T_2614 = _GEN_457 + 4'h1; // @[util.scala 10:8:@5942.6]
  assign _GEN_492 = _T_2614 % 5'h10; // @[util.scala 10:14:@5943.6]
  assign _T_2615 = _GEN_492[4:0]; // @[util.scala 10:14:@5943.6]
  assign _T_2616 = _T_2615 == _GEN_2377; // @[LoadQueue.scala 97:56:@5944.6]
  assign _T_2617 = io_storeEmpty & _T_2616; // @[LoadQueue.scala 96:50:@5945.6]
  assign _T_2619 = _T_2617 == 1'h0; // @[LoadQueue.scala 96:34:@5946.6]
  assign _T_2621 = previousStoreHead <= offsetQ_13; // @[LoadQueue.scala 101:36:@5954.8]
  assign _T_2622 = offsetQ_13 < io_storeHead; // @[LoadQueue.scala 101:86:@5955.8]
  assign _T_2623 = _T_2621 & _T_2622; // @[LoadQueue.scala 101:61:@5956.8]
  assign _T_2626 = io_storeHead <= offsetQ_13; // @[LoadQueue.scala 103:69:@5962.10]
  assign _T_2627 = offsetQ_13 < previousStoreHead; // @[LoadQueue.scala 104:31:@5963.10]
  assign _T_2628 = _T_2626 & _T_2627; // @[LoadQueue.scala 103:94:@5964.10]
  assign _T_2630 = _T_2628 == 1'h0; // @[LoadQueue.scala 103:54:@5965.10]
  assign _T_2631 = _T_2235 & _T_2630; // @[LoadQueue.scala 103:51:@5966.10]
  assign _GEN_820 = _T_2631 ? 1'h0 : checkBits_13; // @[LoadQueue.scala 104:53:@5967.10]
  assign _GEN_821 = _T_2623 ? 1'h0 : _GEN_820; // @[LoadQueue.scala 101:102:@5957.8]
  assign _GEN_822 = io_storeEmpty ? 1'h0 : _GEN_821; // @[LoadQueue.scala 99:27:@5950.6]
  assign _GEN_823 = initBits_13 ? _T_2619 : _GEN_822; // @[LoadQueue.scala 95:34:@5935.4]
  assign _T_2644 = _GEN_491 + 4'h1; // @[util.scala 10:8:@5978.6]
  assign _GEN_510 = _T_2644 % 5'h10; // @[util.scala 10:14:@5979.6]
  assign _T_2645 = _GEN_510[4:0]; // @[util.scala 10:14:@5979.6]
  assign _T_2646 = _T_2645 == _GEN_2377; // @[LoadQueue.scala 97:56:@5980.6]
  assign _T_2647 = io_storeEmpty & _T_2646; // @[LoadQueue.scala 96:50:@5981.6]
  assign _T_2649 = _T_2647 == 1'h0; // @[LoadQueue.scala 96:34:@5982.6]
  assign _T_2651 = previousStoreHead <= offsetQ_14; // @[LoadQueue.scala 101:36:@5990.8]
  assign _T_2652 = offsetQ_14 < io_storeHead; // @[LoadQueue.scala 101:86:@5991.8]
  assign _T_2653 = _T_2651 & _T_2652; // @[LoadQueue.scala 101:61:@5992.8]
  assign _T_2656 = io_storeHead <= offsetQ_14; // @[LoadQueue.scala 103:69:@5998.10]
  assign _T_2657 = offsetQ_14 < previousStoreHead; // @[LoadQueue.scala 104:31:@5999.10]
  assign _T_2658 = _T_2656 & _T_2657; // @[LoadQueue.scala 103:94:@6000.10]
  assign _T_2660 = _T_2658 == 1'h0; // @[LoadQueue.scala 103:54:@6001.10]
  assign _T_2661 = _T_2235 & _T_2660; // @[LoadQueue.scala 103:51:@6002.10]
  assign _GEN_840 = _T_2661 ? 1'h0 : checkBits_14; // @[LoadQueue.scala 104:53:@6003.10]
  assign _GEN_841 = _T_2653 ? 1'h0 : _GEN_840; // @[LoadQueue.scala 101:102:@5993.8]
  assign _GEN_842 = io_storeEmpty ? 1'h0 : _GEN_841; // @[LoadQueue.scala 99:27:@5986.6]
  assign _GEN_843 = initBits_14 ? _T_2649 : _GEN_842; // @[LoadQueue.scala 95:34:@5971.4]
  assign _T_2674 = _GEN_525 + 4'h1; // @[util.scala 10:8:@6014.6]
  assign _GEN_526 = _T_2674 % 5'h10; // @[util.scala 10:14:@6015.6]
  assign _T_2675 = _GEN_526[4:0]; // @[util.scala 10:14:@6015.6]
  assign _T_2676 = _T_2675 == _GEN_2377; // @[LoadQueue.scala 97:56:@6016.6]
  assign _T_2677 = io_storeEmpty & _T_2676; // @[LoadQueue.scala 96:50:@6017.6]
  assign _T_2679 = _T_2677 == 1'h0; // @[LoadQueue.scala 96:34:@6018.6]
  assign _T_2681 = previousStoreHead <= offsetQ_15; // @[LoadQueue.scala 101:36:@6026.8]
  assign _T_2682 = offsetQ_15 < io_storeHead; // @[LoadQueue.scala 101:86:@6027.8]
  assign _T_2683 = _T_2681 & _T_2682; // @[LoadQueue.scala 101:61:@6028.8]
  assign _T_2686 = io_storeHead <= offsetQ_15; // @[LoadQueue.scala 103:69:@6034.10]
  assign _T_2687 = offsetQ_15 < previousStoreHead; // @[LoadQueue.scala 104:31:@6035.10]
  assign _T_2688 = _T_2686 & _T_2687; // @[LoadQueue.scala 103:94:@6036.10]
  assign _T_2690 = _T_2688 == 1'h0; // @[LoadQueue.scala 103:54:@6037.10]
  assign _T_2691 = _T_2235 & _T_2690; // @[LoadQueue.scala 103:51:@6038.10]
  assign _GEN_860 = _T_2691 ? 1'h0 : checkBits_15; // @[LoadQueue.scala 104:53:@6039.10]
  assign _GEN_861 = _T_2683 ? 1'h0 : _GEN_860; // @[LoadQueue.scala 101:102:@6029.8]
  assign _GEN_862 = io_storeEmpty ? 1'h0 : _GEN_861; // @[LoadQueue.scala 99:27:@6022.6]
  assign _GEN_863 = initBits_15 ? _T_2679 : _GEN_862; // @[LoadQueue.scala 95:34:@6007.4]
  assign _T_2695 = 16'h1 << io_storeHead; // @[OneHot.scala 52:12:@6044.4]
  assign _T_2697 = _T_2695[0]; // @[util.scala 60:60:@6046.4]
  assign _T_2698 = _T_2695[1]; // @[util.scala 60:60:@6047.4]
  assign _T_2699 = _T_2695[2]; // @[util.scala 60:60:@6048.4]
  assign _T_2700 = _T_2695[3]; // @[util.scala 60:60:@6049.4]
  assign _T_2701 = _T_2695[4]; // @[util.scala 60:60:@6050.4]
  assign _T_2702 = _T_2695[5]; // @[util.scala 60:60:@6051.4]
  assign _T_2703 = _T_2695[6]; // @[util.scala 60:60:@6052.4]
  assign _T_2704 = _T_2695[7]; // @[util.scala 60:60:@6053.4]
  assign _T_2705 = _T_2695[8]; // @[util.scala 60:60:@6054.4]
  assign _T_2706 = _T_2695[9]; // @[util.scala 60:60:@6055.4]
  assign _T_2707 = _T_2695[10]; // @[util.scala 60:60:@6056.4]
  assign _T_2708 = _T_2695[11]; // @[util.scala 60:60:@6057.4]
  assign _T_2709 = _T_2695[12]; // @[util.scala 60:60:@6058.4]
  assign _T_2710 = _T_2695[13]; // @[util.scala 60:60:@6059.4]
  assign _T_2711 = _T_2695[14]; // @[util.scala 60:60:@6060.4]
  assign _T_2712 = _T_2695[15]; // @[util.scala 60:60:@6061.4]
  assign _T_4843 = {io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0}; // @[Mux.scala 19:72:@7585.4]
  assign _T_4850 = {io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8}; // @[Mux.scala 19:72:@7592.4]
  assign _T_4851 = {io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,_T_4843}; // @[Mux.scala 19:72:@7593.4]
  assign _T_4853 = _T_2697 ? _T_4851 : 512'h0; // @[Mux.scala 19:72:@7594.4]
  assign _T_4860 = {io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1}; // @[Mux.scala 19:72:@7601.4]
  assign _T_4867 = {io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9}; // @[Mux.scala 19:72:@7608.4]
  assign _T_4868 = {io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,_T_4860}; // @[Mux.scala 19:72:@7609.4]
  assign _T_4870 = _T_2698 ? _T_4868 : 512'h0; // @[Mux.scala 19:72:@7610.4]
  assign _T_4877 = {io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2}; // @[Mux.scala 19:72:@7617.4]
  assign _T_4884 = {io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10}; // @[Mux.scala 19:72:@7624.4]
  assign _T_4885 = {io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,_T_4877}; // @[Mux.scala 19:72:@7625.4]
  assign _T_4887 = _T_2699 ? _T_4885 : 512'h0; // @[Mux.scala 19:72:@7626.4]
  assign _T_4894 = {io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3}; // @[Mux.scala 19:72:@7633.4]
  assign _T_4901 = {io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11}; // @[Mux.scala 19:72:@7640.4]
  assign _T_4902 = {io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,_T_4894}; // @[Mux.scala 19:72:@7641.4]
  assign _T_4904 = _T_2700 ? _T_4902 : 512'h0; // @[Mux.scala 19:72:@7642.4]
  assign _T_4911 = {io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4}; // @[Mux.scala 19:72:@7649.4]
  assign _T_4918 = {io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12}; // @[Mux.scala 19:72:@7656.4]
  assign _T_4919 = {io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,_T_4911}; // @[Mux.scala 19:72:@7657.4]
  assign _T_4921 = _T_2701 ? _T_4919 : 512'h0; // @[Mux.scala 19:72:@7658.4]
  assign _T_4928 = {io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5}; // @[Mux.scala 19:72:@7665.4]
  assign _T_4935 = {io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13}; // @[Mux.scala 19:72:@7672.4]
  assign _T_4936 = {io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,_T_4928}; // @[Mux.scala 19:72:@7673.4]
  assign _T_4938 = _T_2702 ? _T_4936 : 512'h0; // @[Mux.scala 19:72:@7674.4]
  assign _T_4945 = {io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6}; // @[Mux.scala 19:72:@7681.4]
  assign _T_4952 = {io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14}; // @[Mux.scala 19:72:@7688.4]
  assign _T_4953 = {io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,_T_4945}; // @[Mux.scala 19:72:@7689.4]
  assign _T_4955 = _T_2703 ? _T_4953 : 512'h0; // @[Mux.scala 19:72:@7690.4]
  assign _T_4962 = {io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7}; // @[Mux.scala 19:72:@7697.4]
  assign _T_4969 = {io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15}; // @[Mux.scala 19:72:@7704.4]
  assign _T_4970 = {io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,_T_4962}; // @[Mux.scala 19:72:@7705.4]
  assign _T_4972 = _T_2704 ? _T_4970 : 512'h0; // @[Mux.scala 19:72:@7706.4]
  assign _T_4987 = {io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,_T_4850}; // @[Mux.scala 19:72:@7721.4]
  assign _T_4989 = _T_2705 ? _T_4987 : 512'h0; // @[Mux.scala 19:72:@7722.4]
  assign _T_5004 = {io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,_T_4867}; // @[Mux.scala 19:72:@7737.4]
  assign _T_5006 = _T_2706 ? _T_5004 : 512'h0; // @[Mux.scala 19:72:@7738.4]
  assign _T_5021 = {io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,_T_4884}; // @[Mux.scala 19:72:@7753.4]
  assign _T_5023 = _T_2707 ? _T_5021 : 512'h0; // @[Mux.scala 19:72:@7754.4]
  assign _T_5038 = {io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,_T_4901}; // @[Mux.scala 19:72:@7769.4]
  assign _T_5040 = _T_2708 ? _T_5038 : 512'h0; // @[Mux.scala 19:72:@7770.4]
  assign _T_5055 = {io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,_T_4918}; // @[Mux.scala 19:72:@7785.4]
  assign _T_5057 = _T_2709 ? _T_5055 : 512'h0; // @[Mux.scala 19:72:@7786.4]
  assign _T_5072 = {io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,_T_4935}; // @[Mux.scala 19:72:@7801.4]
  assign _T_5074 = _T_2710 ? _T_5072 : 512'h0; // @[Mux.scala 19:72:@7802.4]
  assign _T_5089 = {io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,_T_4952}; // @[Mux.scala 19:72:@7817.4]
  assign _T_5091 = _T_2711 ? _T_5089 : 512'h0; // @[Mux.scala 19:72:@7818.4]
  assign _T_5106 = {io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,_T_4969}; // @[Mux.scala 19:72:@7833.4]
  assign _T_5108 = _T_2712 ? _T_5106 : 512'h0; // @[Mux.scala 19:72:@7834.4]
  assign _T_5109 = _T_4853 | _T_4870; // @[Mux.scala 19:72:@7835.4]
  assign _T_5110 = _T_5109 | _T_4887; // @[Mux.scala 19:72:@7836.4]
  assign _T_5111 = _T_5110 | _T_4904; // @[Mux.scala 19:72:@7837.4]
  assign _T_5112 = _T_5111 | _T_4921; // @[Mux.scala 19:72:@7838.4]
  assign _T_5113 = _T_5112 | _T_4938; // @[Mux.scala 19:72:@7839.4]
  assign _T_5114 = _T_5113 | _T_4955; // @[Mux.scala 19:72:@7840.4]
  assign _T_5115 = _T_5114 | _T_4972; // @[Mux.scala 19:72:@7841.4]
  assign _T_5116 = _T_5115 | _T_4989; // @[Mux.scala 19:72:@7842.4]
  assign _T_5117 = _T_5116 | _T_5006; // @[Mux.scala 19:72:@7843.4]
  assign _T_5118 = _T_5117 | _T_5023; // @[Mux.scala 19:72:@7844.4]
  assign _T_5119 = _T_5118 | _T_5040; // @[Mux.scala 19:72:@7845.4]
  assign _T_5120 = _T_5119 | _T_5057; // @[Mux.scala 19:72:@7846.4]
  assign _T_5121 = _T_5120 | _T_5074; // @[Mux.scala 19:72:@7847.4]
  assign _T_5122 = _T_5121 | _T_5091; // @[Mux.scala 19:72:@7848.4]
  assign _T_5123 = _T_5122 | _T_5108; // @[Mux.scala 19:72:@7849.4]
  assign _T_5700 = {io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0}; // @[Mux.scala 19:72:@8199.4]
  assign _T_5707 = {io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8}; // @[Mux.scala 19:72:@8206.4]
  assign _T_5708 = {io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,_T_5700}; // @[Mux.scala 19:72:@8207.4]
  assign _T_5710 = _T_2697 ? _T_5708 : 16'h0; // @[Mux.scala 19:72:@8208.4]
  assign _T_5717 = {io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1}; // @[Mux.scala 19:72:@8215.4]
  assign _T_5724 = {io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9}; // @[Mux.scala 19:72:@8222.4]
  assign _T_5725 = {io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,_T_5717}; // @[Mux.scala 19:72:@8223.4]
  assign _T_5727 = _T_2698 ? _T_5725 : 16'h0; // @[Mux.scala 19:72:@8224.4]
  assign _T_5734 = {io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2}; // @[Mux.scala 19:72:@8231.4]
  assign _T_5741 = {io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10}; // @[Mux.scala 19:72:@8238.4]
  assign _T_5742 = {io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,_T_5734}; // @[Mux.scala 19:72:@8239.4]
  assign _T_5744 = _T_2699 ? _T_5742 : 16'h0; // @[Mux.scala 19:72:@8240.4]
  assign _T_5751 = {io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3}; // @[Mux.scala 19:72:@8247.4]
  assign _T_5758 = {io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11}; // @[Mux.scala 19:72:@8254.4]
  assign _T_5759 = {io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,_T_5751}; // @[Mux.scala 19:72:@8255.4]
  assign _T_5761 = _T_2700 ? _T_5759 : 16'h0; // @[Mux.scala 19:72:@8256.4]
  assign _T_5768 = {io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4}; // @[Mux.scala 19:72:@8263.4]
  assign _T_5775 = {io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12}; // @[Mux.scala 19:72:@8270.4]
  assign _T_5776 = {io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,_T_5768}; // @[Mux.scala 19:72:@8271.4]
  assign _T_5778 = _T_2701 ? _T_5776 : 16'h0; // @[Mux.scala 19:72:@8272.4]
  assign _T_5785 = {io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5}; // @[Mux.scala 19:72:@8279.4]
  assign _T_5792 = {io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13}; // @[Mux.scala 19:72:@8286.4]
  assign _T_5793 = {io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,_T_5785}; // @[Mux.scala 19:72:@8287.4]
  assign _T_5795 = _T_2702 ? _T_5793 : 16'h0; // @[Mux.scala 19:72:@8288.4]
  assign _T_5802 = {io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6}; // @[Mux.scala 19:72:@8295.4]
  assign _T_5809 = {io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14}; // @[Mux.scala 19:72:@8302.4]
  assign _T_5810 = {io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,_T_5802}; // @[Mux.scala 19:72:@8303.4]
  assign _T_5812 = _T_2703 ? _T_5810 : 16'h0; // @[Mux.scala 19:72:@8304.4]
  assign _T_5819 = {io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7}; // @[Mux.scala 19:72:@8311.4]
  assign _T_5826 = {io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15}; // @[Mux.scala 19:72:@8318.4]
  assign _T_5827 = {io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,_T_5819}; // @[Mux.scala 19:72:@8319.4]
  assign _T_5829 = _T_2704 ? _T_5827 : 16'h0; // @[Mux.scala 19:72:@8320.4]
  assign _T_5844 = {io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,_T_5707}; // @[Mux.scala 19:72:@8335.4]
  assign _T_5846 = _T_2705 ? _T_5844 : 16'h0; // @[Mux.scala 19:72:@8336.4]
  assign _T_5861 = {io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,_T_5724}; // @[Mux.scala 19:72:@8351.4]
  assign _T_5863 = _T_2706 ? _T_5861 : 16'h0; // @[Mux.scala 19:72:@8352.4]
  assign _T_5878 = {io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,_T_5741}; // @[Mux.scala 19:72:@8367.4]
  assign _T_5880 = _T_2707 ? _T_5878 : 16'h0; // @[Mux.scala 19:72:@8368.4]
  assign _T_5895 = {io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,_T_5758}; // @[Mux.scala 19:72:@8383.4]
  assign _T_5897 = _T_2708 ? _T_5895 : 16'h0; // @[Mux.scala 19:72:@8384.4]
  assign _T_5912 = {io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,_T_5775}; // @[Mux.scala 19:72:@8399.4]
  assign _T_5914 = _T_2709 ? _T_5912 : 16'h0; // @[Mux.scala 19:72:@8400.4]
  assign _T_5929 = {io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,_T_5792}; // @[Mux.scala 19:72:@8415.4]
  assign _T_5931 = _T_2710 ? _T_5929 : 16'h0; // @[Mux.scala 19:72:@8416.4]
  assign _T_5946 = {io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,_T_5809}; // @[Mux.scala 19:72:@8431.4]
  assign _T_5948 = _T_2711 ? _T_5946 : 16'h0; // @[Mux.scala 19:72:@8432.4]
  assign _T_5963 = {io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,_T_5826}; // @[Mux.scala 19:72:@8447.4]
  assign _T_5965 = _T_2712 ? _T_5963 : 16'h0; // @[Mux.scala 19:72:@8448.4]
  assign _T_5966 = _T_5710 | _T_5727; // @[Mux.scala 19:72:@8449.4]
  assign _T_5967 = _T_5966 | _T_5744; // @[Mux.scala 19:72:@8450.4]
  assign _T_5968 = _T_5967 | _T_5761; // @[Mux.scala 19:72:@8451.4]
  assign _T_5969 = _T_5968 | _T_5778; // @[Mux.scala 19:72:@8452.4]
  assign _T_5970 = _T_5969 | _T_5795; // @[Mux.scala 19:72:@8453.4]
  assign _T_5971 = _T_5970 | _T_5812; // @[Mux.scala 19:72:@8454.4]
  assign _T_5972 = _T_5971 | _T_5829; // @[Mux.scala 19:72:@8455.4]
  assign _T_5973 = _T_5972 | _T_5846; // @[Mux.scala 19:72:@8456.4]
  assign _T_5974 = _T_5973 | _T_5863; // @[Mux.scala 19:72:@8457.4]
  assign _T_5975 = _T_5974 | _T_5880; // @[Mux.scala 19:72:@8458.4]
  assign _T_5976 = _T_5975 | _T_5897; // @[Mux.scala 19:72:@8459.4]
  assign _T_5977 = _T_5976 | _T_5914; // @[Mux.scala 19:72:@8460.4]
  assign _T_5978 = _T_5977 | _T_5931; // @[Mux.scala 19:72:@8461.4]
  assign _T_5979 = _T_5978 | _T_5948; // @[Mux.scala 19:72:@8462.4]
  assign _T_5980 = _T_5979 | _T_5965; // @[Mux.scala 19:72:@8463.4]
  assign _T_6121 = io_storeHead < io_storeTail; // @[LoadQueue.scala 121:105:@8499.4]
  assign _T_6123 = io_storeHead <= 4'h0; // @[LoadQueue.scala 122:18:@8500.4]
  assign _T_6125 = 4'h0 < io_storeTail; // @[LoadQueue.scala 122:36:@8501.4]
  assign _T_6126 = _T_6123 & _T_6125; // @[LoadQueue.scala 122:27:@8502.4]
  assign _T_6128 = io_storeEmpty == 1'h0; // @[LoadQueue.scala 122:52:@8503.4]
  assign _T_6130 = io_storeTail <= 4'h0; // @[LoadQueue.scala 122:85:@8504.4]
  assign _T_6132 = 4'h0 < io_storeHead; // @[LoadQueue.scala 122:103:@8505.4]
  assign _T_6133 = _T_6130 & _T_6132; // @[LoadQueue.scala 122:94:@8506.4]
  assign _T_6135 = _T_6133 == 1'h0; // @[LoadQueue.scala 122:70:@8507.4]
  assign _T_6136 = _T_6128 & _T_6135; // @[LoadQueue.scala 122:67:@8508.4]
  assign validEntriesInStoreQ_0 = _T_6121 ? _T_6126 : _T_6136; // @[LoadQueue.scala 121:91:@8509.4]
  assign _T_6140 = io_storeHead <= 4'h1; // @[LoadQueue.scala 122:18:@8511.4]
  assign _T_6142 = 4'h1 < io_storeTail; // @[LoadQueue.scala 122:36:@8512.4]
  assign _T_6143 = _T_6140 & _T_6142; // @[LoadQueue.scala 122:27:@8513.4]
  assign _T_6147 = io_storeTail <= 4'h1; // @[LoadQueue.scala 122:85:@8515.4]
  assign _T_6149 = 4'h1 < io_storeHead; // @[LoadQueue.scala 122:103:@8516.4]
  assign _T_6150 = _T_6147 & _T_6149; // @[LoadQueue.scala 122:94:@8517.4]
  assign _T_6152 = _T_6150 == 1'h0; // @[LoadQueue.scala 122:70:@8518.4]
  assign _T_6153 = _T_6128 & _T_6152; // @[LoadQueue.scala 122:67:@8519.4]
  assign validEntriesInStoreQ_1 = _T_6121 ? _T_6143 : _T_6153; // @[LoadQueue.scala 121:91:@8520.4]
  assign _T_6157 = io_storeHead <= 4'h2; // @[LoadQueue.scala 122:18:@8522.4]
  assign _T_6159 = 4'h2 < io_storeTail; // @[LoadQueue.scala 122:36:@8523.4]
  assign _T_6160 = _T_6157 & _T_6159; // @[LoadQueue.scala 122:27:@8524.4]
  assign _T_6164 = io_storeTail <= 4'h2; // @[LoadQueue.scala 122:85:@8526.4]
  assign _T_6166 = 4'h2 < io_storeHead; // @[LoadQueue.scala 122:103:@8527.4]
  assign _T_6167 = _T_6164 & _T_6166; // @[LoadQueue.scala 122:94:@8528.4]
  assign _T_6169 = _T_6167 == 1'h0; // @[LoadQueue.scala 122:70:@8529.4]
  assign _T_6170 = _T_6128 & _T_6169; // @[LoadQueue.scala 122:67:@8530.4]
  assign validEntriesInStoreQ_2 = _T_6121 ? _T_6160 : _T_6170; // @[LoadQueue.scala 121:91:@8531.4]
  assign _T_6174 = io_storeHead <= 4'h3; // @[LoadQueue.scala 122:18:@8533.4]
  assign _T_6176 = 4'h3 < io_storeTail; // @[LoadQueue.scala 122:36:@8534.4]
  assign _T_6177 = _T_6174 & _T_6176; // @[LoadQueue.scala 122:27:@8535.4]
  assign _T_6181 = io_storeTail <= 4'h3; // @[LoadQueue.scala 122:85:@8537.4]
  assign _T_6183 = 4'h3 < io_storeHead; // @[LoadQueue.scala 122:103:@8538.4]
  assign _T_6184 = _T_6181 & _T_6183; // @[LoadQueue.scala 122:94:@8539.4]
  assign _T_6186 = _T_6184 == 1'h0; // @[LoadQueue.scala 122:70:@8540.4]
  assign _T_6187 = _T_6128 & _T_6186; // @[LoadQueue.scala 122:67:@8541.4]
  assign validEntriesInStoreQ_3 = _T_6121 ? _T_6177 : _T_6187; // @[LoadQueue.scala 121:91:@8542.4]
  assign _T_6191 = io_storeHead <= 4'h4; // @[LoadQueue.scala 122:18:@8544.4]
  assign _T_6193 = 4'h4 < io_storeTail; // @[LoadQueue.scala 122:36:@8545.4]
  assign _T_6194 = _T_6191 & _T_6193; // @[LoadQueue.scala 122:27:@8546.4]
  assign _T_6198 = io_storeTail <= 4'h4; // @[LoadQueue.scala 122:85:@8548.4]
  assign _T_6200 = 4'h4 < io_storeHead; // @[LoadQueue.scala 122:103:@8549.4]
  assign _T_6201 = _T_6198 & _T_6200; // @[LoadQueue.scala 122:94:@8550.4]
  assign _T_6203 = _T_6201 == 1'h0; // @[LoadQueue.scala 122:70:@8551.4]
  assign _T_6204 = _T_6128 & _T_6203; // @[LoadQueue.scala 122:67:@8552.4]
  assign validEntriesInStoreQ_4 = _T_6121 ? _T_6194 : _T_6204; // @[LoadQueue.scala 121:91:@8553.4]
  assign _T_6208 = io_storeHead <= 4'h5; // @[LoadQueue.scala 122:18:@8555.4]
  assign _T_6210 = 4'h5 < io_storeTail; // @[LoadQueue.scala 122:36:@8556.4]
  assign _T_6211 = _T_6208 & _T_6210; // @[LoadQueue.scala 122:27:@8557.4]
  assign _T_6215 = io_storeTail <= 4'h5; // @[LoadQueue.scala 122:85:@8559.4]
  assign _T_6217 = 4'h5 < io_storeHead; // @[LoadQueue.scala 122:103:@8560.4]
  assign _T_6218 = _T_6215 & _T_6217; // @[LoadQueue.scala 122:94:@8561.4]
  assign _T_6220 = _T_6218 == 1'h0; // @[LoadQueue.scala 122:70:@8562.4]
  assign _T_6221 = _T_6128 & _T_6220; // @[LoadQueue.scala 122:67:@8563.4]
  assign validEntriesInStoreQ_5 = _T_6121 ? _T_6211 : _T_6221; // @[LoadQueue.scala 121:91:@8564.4]
  assign _T_6225 = io_storeHead <= 4'h6; // @[LoadQueue.scala 122:18:@8566.4]
  assign _T_6227 = 4'h6 < io_storeTail; // @[LoadQueue.scala 122:36:@8567.4]
  assign _T_6228 = _T_6225 & _T_6227; // @[LoadQueue.scala 122:27:@8568.4]
  assign _T_6232 = io_storeTail <= 4'h6; // @[LoadQueue.scala 122:85:@8570.4]
  assign _T_6234 = 4'h6 < io_storeHead; // @[LoadQueue.scala 122:103:@8571.4]
  assign _T_6235 = _T_6232 & _T_6234; // @[LoadQueue.scala 122:94:@8572.4]
  assign _T_6237 = _T_6235 == 1'h0; // @[LoadQueue.scala 122:70:@8573.4]
  assign _T_6238 = _T_6128 & _T_6237; // @[LoadQueue.scala 122:67:@8574.4]
  assign validEntriesInStoreQ_6 = _T_6121 ? _T_6228 : _T_6238; // @[LoadQueue.scala 121:91:@8575.4]
  assign _T_6242 = io_storeHead <= 4'h7; // @[LoadQueue.scala 122:18:@8577.4]
  assign _T_6244 = 4'h7 < io_storeTail; // @[LoadQueue.scala 122:36:@8578.4]
  assign _T_6245 = _T_6242 & _T_6244; // @[LoadQueue.scala 122:27:@8579.4]
  assign _T_6249 = io_storeTail <= 4'h7; // @[LoadQueue.scala 122:85:@8581.4]
  assign _T_6251 = 4'h7 < io_storeHead; // @[LoadQueue.scala 122:103:@8582.4]
  assign _T_6252 = _T_6249 & _T_6251; // @[LoadQueue.scala 122:94:@8583.4]
  assign _T_6254 = _T_6252 == 1'h0; // @[LoadQueue.scala 122:70:@8584.4]
  assign _T_6255 = _T_6128 & _T_6254; // @[LoadQueue.scala 122:67:@8585.4]
  assign validEntriesInStoreQ_7 = _T_6121 ? _T_6245 : _T_6255; // @[LoadQueue.scala 121:91:@8586.4]
  assign _T_6259 = io_storeHead <= 4'h8; // @[LoadQueue.scala 122:18:@8588.4]
  assign _T_6261 = 4'h8 < io_storeTail; // @[LoadQueue.scala 122:36:@8589.4]
  assign _T_6262 = _T_6259 & _T_6261; // @[LoadQueue.scala 122:27:@8590.4]
  assign _T_6266 = io_storeTail <= 4'h8; // @[LoadQueue.scala 122:85:@8592.4]
  assign _T_6268 = 4'h8 < io_storeHead; // @[LoadQueue.scala 122:103:@8593.4]
  assign _T_6269 = _T_6266 & _T_6268; // @[LoadQueue.scala 122:94:@8594.4]
  assign _T_6271 = _T_6269 == 1'h0; // @[LoadQueue.scala 122:70:@8595.4]
  assign _T_6272 = _T_6128 & _T_6271; // @[LoadQueue.scala 122:67:@8596.4]
  assign validEntriesInStoreQ_8 = _T_6121 ? _T_6262 : _T_6272; // @[LoadQueue.scala 121:91:@8597.4]
  assign _T_6276 = io_storeHead <= 4'h9; // @[LoadQueue.scala 122:18:@8599.4]
  assign _T_6278 = 4'h9 < io_storeTail; // @[LoadQueue.scala 122:36:@8600.4]
  assign _T_6279 = _T_6276 & _T_6278; // @[LoadQueue.scala 122:27:@8601.4]
  assign _T_6283 = io_storeTail <= 4'h9; // @[LoadQueue.scala 122:85:@8603.4]
  assign _T_6285 = 4'h9 < io_storeHead; // @[LoadQueue.scala 122:103:@8604.4]
  assign _T_6286 = _T_6283 & _T_6285; // @[LoadQueue.scala 122:94:@8605.4]
  assign _T_6288 = _T_6286 == 1'h0; // @[LoadQueue.scala 122:70:@8606.4]
  assign _T_6289 = _T_6128 & _T_6288; // @[LoadQueue.scala 122:67:@8607.4]
  assign validEntriesInStoreQ_9 = _T_6121 ? _T_6279 : _T_6289; // @[LoadQueue.scala 121:91:@8608.4]
  assign _T_6293 = io_storeHead <= 4'ha; // @[LoadQueue.scala 122:18:@8610.4]
  assign _T_6295 = 4'ha < io_storeTail; // @[LoadQueue.scala 122:36:@8611.4]
  assign _T_6296 = _T_6293 & _T_6295; // @[LoadQueue.scala 122:27:@8612.4]
  assign _T_6300 = io_storeTail <= 4'ha; // @[LoadQueue.scala 122:85:@8614.4]
  assign _T_6302 = 4'ha < io_storeHead; // @[LoadQueue.scala 122:103:@8615.4]
  assign _T_6303 = _T_6300 & _T_6302; // @[LoadQueue.scala 122:94:@8616.4]
  assign _T_6305 = _T_6303 == 1'h0; // @[LoadQueue.scala 122:70:@8617.4]
  assign _T_6306 = _T_6128 & _T_6305; // @[LoadQueue.scala 122:67:@8618.4]
  assign validEntriesInStoreQ_10 = _T_6121 ? _T_6296 : _T_6306; // @[LoadQueue.scala 121:91:@8619.4]
  assign _T_6310 = io_storeHead <= 4'hb; // @[LoadQueue.scala 122:18:@8621.4]
  assign _T_6312 = 4'hb < io_storeTail; // @[LoadQueue.scala 122:36:@8622.4]
  assign _T_6313 = _T_6310 & _T_6312; // @[LoadQueue.scala 122:27:@8623.4]
  assign _T_6317 = io_storeTail <= 4'hb; // @[LoadQueue.scala 122:85:@8625.4]
  assign _T_6319 = 4'hb < io_storeHead; // @[LoadQueue.scala 122:103:@8626.4]
  assign _T_6320 = _T_6317 & _T_6319; // @[LoadQueue.scala 122:94:@8627.4]
  assign _T_6322 = _T_6320 == 1'h0; // @[LoadQueue.scala 122:70:@8628.4]
  assign _T_6323 = _T_6128 & _T_6322; // @[LoadQueue.scala 122:67:@8629.4]
  assign validEntriesInStoreQ_11 = _T_6121 ? _T_6313 : _T_6323; // @[LoadQueue.scala 121:91:@8630.4]
  assign _T_6327 = io_storeHead <= 4'hc; // @[LoadQueue.scala 122:18:@8632.4]
  assign _T_6329 = 4'hc < io_storeTail; // @[LoadQueue.scala 122:36:@8633.4]
  assign _T_6330 = _T_6327 & _T_6329; // @[LoadQueue.scala 122:27:@8634.4]
  assign _T_6334 = io_storeTail <= 4'hc; // @[LoadQueue.scala 122:85:@8636.4]
  assign _T_6336 = 4'hc < io_storeHead; // @[LoadQueue.scala 122:103:@8637.4]
  assign _T_6337 = _T_6334 & _T_6336; // @[LoadQueue.scala 122:94:@8638.4]
  assign _T_6339 = _T_6337 == 1'h0; // @[LoadQueue.scala 122:70:@8639.4]
  assign _T_6340 = _T_6128 & _T_6339; // @[LoadQueue.scala 122:67:@8640.4]
  assign validEntriesInStoreQ_12 = _T_6121 ? _T_6330 : _T_6340; // @[LoadQueue.scala 121:91:@8641.4]
  assign _T_6344 = io_storeHead <= 4'hd; // @[LoadQueue.scala 122:18:@8643.4]
  assign _T_6346 = 4'hd < io_storeTail; // @[LoadQueue.scala 122:36:@8644.4]
  assign _T_6347 = _T_6344 & _T_6346; // @[LoadQueue.scala 122:27:@8645.4]
  assign _T_6351 = io_storeTail <= 4'hd; // @[LoadQueue.scala 122:85:@8647.4]
  assign _T_6353 = 4'hd < io_storeHead; // @[LoadQueue.scala 122:103:@8648.4]
  assign _T_6354 = _T_6351 & _T_6353; // @[LoadQueue.scala 122:94:@8649.4]
  assign _T_6356 = _T_6354 == 1'h0; // @[LoadQueue.scala 122:70:@8650.4]
  assign _T_6357 = _T_6128 & _T_6356; // @[LoadQueue.scala 122:67:@8651.4]
  assign validEntriesInStoreQ_13 = _T_6121 ? _T_6347 : _T_6357; // @[LoadQueue.scala 121:91:@8652.4]
  assign _T_6361 = io_storeHead <= 4'he; // @[LoadQueue.scala 122:18:@8654.4]
  assign _T_6363 = 4'he < io_storeTail; // @[LoadQueue.scala 122:36:@8655.4]
  assign _T_6364 = _T_6361 & _T_6363; // @[LoadQueue.scala 122:27:@8656.4]
  assign _T_6368 = io_storeTail <= 4'he; // @[LoadQueue.scala 122:85:@8658.4]
  assign _T_6370 = 4'he < io_storeHead; // @[LoadQueue.scala 122:103:@8659.4]
  assign _T_6371 = _T_6368 & _T_6370; // @[LoadQueue.scala 122:94:@8660.4]
  assign _T_6373 = _T_6371 == 1'h0; // @[LoadQueue.scala 122:70:@8661.4]
  assign _T_6374 = _T_6128 & _T_6373; // @[LoadQueue.scala 122:67:@8662.4]
  assign validEntriesInStoreQ_14 = _T_6121 ? _T_6364 : _T_6374; // @[LoadQueue.scala 121:91:@8663.4]
  assign validEntriesInStoreQ_15 = _T_6121 ? 1'h0 : _T_6128; // @[LoadQueue.scala 121:91:@8674.4]
  assign storesToCheck_0_0 = _T_2236 ? _T_6123 : 1'h1; // @[LoadQueue.scala 131:10:@8701.4]
  assign _T_7662 = 4'h1 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8704.4]
  assign _T_7663 = _T_6140 & _T_7662; // @[LoadQueue.scala 131:72:@8705.4]
  assign _T_7665 = offsetQ_0 < 4'h1; // @[LoadQueue.scala 132:33:@8706.4]
  assign _T_7668 = _T_7665 & _T_6149; // @[LoadQueue.scala 132:41:@8708.4]
  assign _T_7670 = _T_7668 == 1'h0; // @[LoadQueue.scala 132:9:@8709.4]
  assign storesToCheck_0_1 = _T_2236 ? _T_7663 : _T_7670; // @[LoadQueue.scala 131:10:@8710.4]
  assign _T_7676 = 4'h2 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8713.4]
  assign _T_7677 = _T_6157 & _T_7676; // @[LoadQueue.scala 131:72:@8714.4]
  assign _T_7679 = offsetQ_0 < 4'h2; // @[LoadQueue.scala 132:33:@8715.4]
  assign _T_7682 = _T_7679 & _T_6166; // @[LoadQueue.scala 132:41:@8717.4]
  assign _T_7684 = _T_7682 == 1'h0; // @[LoadQueue.scala 132:9:@8718.4]
  assign storesToCheck_0_2 = _T_2236 ? _T_7677 : _T_7684; // @[LoadQueue.scala 131:10:@8719.4]
  assign _T_7690 = 4'h3 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8722.4]
  assign _T_7691 = _T_6174 & _T_7690; // @[LoadQueue.scala 131:72:@8723.4]
  assign _T_7693 = offsetQ_0 < 4'h3; // @[LoadQueue.scala 132:33:@8724.4]
  assign _T_7696 = _T_7693 & _T_6183; // @[LoadQueue.scala 132:41:@8726.4]
  assign _T_7698 = _T_7696 == 1'h0; // @[LoadQueue.scala 132:9:@8727.4]
  assign storesToCheck_0_3 = _T_2236 ? _T_7691 : _T_7698; // @[LoadQueue.scala 131:10:@8728.4]
  assign _T_7704 = 4'h4 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8731.4]
  assign _T_7705 = _T_6191 & _T_7704; // @[LoadQueue.scala 131:72:@8732.4]
  assign _T_7707 = offsetQ_0 < 4'h4; // @[LoadQueue.scala 132:33:@8733.4]
  assign _T_7710 = _T_7707 & _T_6200; // @[LoadQueue.scala 132:41:@8735.4]
  assign _T_7712 = _T_7710 == 1'h0; // @[LoadQueue.scala 132:9:@8736.4]
  assign storesToCheck_0_4 = _T_2236 ? _T_7705 : _T_7712; // @[LoadQueue.scala 131:10:@8737.4]
  assign _T_7718 = 4'h5 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8740.4]
  assign _T_7719 = _T_6208 & _T_7718; // @[LoadQueue.scala 131:72:@8741.4]
  assign _T_7721 = offsetQ_0 < 4'h5; // @[LoadQueue.scala 132:33:@8742.4]
  assign _T_7724 = _T_7721 & _T_6217; // @[LoadQueue.scala 132:41:@8744.4]
  assign _T_7726 = _T_7724 == 1'h0; // @[LoadQueue.scala 132:9:@8745.4]
  assign storesToCheck_0_5 = _T_2236 ? _T_7719 : _T_7726; // @[LoadQueue.scala 131:10:@8746.4]
  assign _T_7732 = 4'h6 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8749.4]
  assign _T_7733 = _T_6225 & _T_7732; // @[LoadQueue.scala 131:72:@8750.4]
  assign _T_7735 = offsetQ_0 < 4'h6; // @[LoadQueue.scala 132:33:@8751.4]
  assign _T_7738 = _T_7735 & _T_6234; // @[LoadQueue.scala 132:41:@8753.4]
  assign _T_7740 = _T_7738 == 1'h0; // @[LoadQueue.scala 132:9:@8754.4]
  assign storesToCheck_0_6 = _T_2236 ? _T_7733 : _T_7740; // @[LoadQueue.scala 131:10:@8755.4]
  assign _T_7746 = 4'h7 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8758.4]
  assign _T_7747 = _T_6242 & _T_7746; // @[LoadQueue.scala 131:72:@8759.4]
  assign _T_7749 = offsetQ_0 < 4'h7; // @[LoadQueue.scala 132:33:@8760.4]
  assign _T_7752 = _T_7749 & _T_6251; // @[LoadQueue.scala 132:41:@8762.4]
  assign _T_7754 = _T_7752 == 1'h0; // @[LoadQueue.scala 132:9:@8763.4]
  assign storesToCheck_0_7 = _T_2236 ? _T_7747 : _T_7754; // @[LoadQueue.scala 131:10:@8764.4]
  assign _T_7760 = 4'h8 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8767.4]
  assign _T_7761 = _T_6259 & _T_7760; // @[LoadQueue.scala 131:72:@8768.4]
  assign _T_7763 = offsetQ_0 < 4'h8; // @[LoadQueue.scala 132:33:@8769.4]
  assign _T_7766 = _T_7763 & _T_6268; // @[LoadQueue.scala 132:41:@8771.4]
  assign _T_7768 = _T_7766 == 1'h0; // @[LoadQueue.scala 132:9:@8772.4]
  assign storesToCheck_0_8 = _T_2236 ? _T_7761 : _T_7768; // @[LoadQueue.scala 131:10:@8773.4]
  assign _T_7774 = 4'h9 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8776.4]
  assign _T_7775 = _T_6276 & _T_7774; // @[LoadQueue.scala 131:72:@8777.4]
  assign _T_7777 = offsetQ_0 < 4'h9; // @[LoadQueue.scala 132:33:@8778.4]
  assign _T_7780 = _T_7777 & _T_6285; // @[LoadQueue.scala 132:41:@8780.4]
  assign _T_7782 = _T_7780 == 1'h0; // @[LoadQueue.scala 132:9:@8781.4]
  assign storesToCheck_0_9 = _T_2236 ? _T_7775 : _T_7782; // @[LoadQueue.scala 131:10:@8782.4]
  assign _T_7788 = 4'ha <= offsetQ_0; // @[LoadQueue.scala 131:81:@8785.4]
  assign _T_7789 = _T_6293 & _T_7788; // @[LoadQueue.scala 131:72:@8786.4]
  assign _T_7791 = offsetQ_0 < 4'ha; // @[LoadQueue.scala 132:33:@8787.4]
  assign _T_7794 = _T_7791 & _T_6302; // @[LoadQueue.scala 132:41:@8789.4]
  assign _T_7796 = _T_7794 == 1'h0; // @[LoadQueue.scala 132:9:@8790.4]
  assign storesToCheck_0_10 = _T_2236 ? _T_7789 : _T_7796; // @[LoadQueue.scala 131:10:@8791.4]
  assign _T_7802 = 4'hb <= offsetQ_0; // @[LoadQueue.scala 131:81:@8794.4]
  assign _T_7803 = _T_6310 & _T_7802; // @[LoadQueue.scala 131:72:@8795.4]
  assign _T_7805 = offsetQ_0 < 4'hb; // @[LoadQueue.scala 132:33:@8796.4]
  assign _T_7808 = _T_7805 & _T_6319; // @[LoadQueue.scala 132:41:@8798.4]
  assign _T_7810 = _T_7808 == 1'h0; // @[LoadQueue.scala 132:9:@8799.4]
  assign storesToCheck_0_11 = _T_2236 ? _T_7803 : _T_7810; // @[LoadQueue.scala 131:10:@8800.4]
  assign _T_7816 = 4'hc <= offsetQ_0; // @[LoadQueue.scala 131:81:@8803.4]
  assign _T_7817 = _T_6327 & _T_7816; // @[LoadQueue.scala 131:72:@8804.4]
  assign _T_7819 = offsetQ_0 < 4'hc; // @[LoadQueue.scala 132:33:@8805.4]
  assign _T_7822 = _T_7819 & _T_6336; // @[LoadQueue.scala 132:41:@8807.4]
  assign _T_7824 = _T_7822 == 1'h0; // @[LoadQueue.scala 132:9:@8808.4]
  assign storesToCheck_0_12 = _T_2236 ? _T_7817 : _T_7824; // @[LoadQueue.scala 131:10:@8809.4]
  assign _T_7830 = 4'hd <= offsetQ_0; // @[LoadQueue.scala 131:81:@8812.4]
  assign _T_7831 = _T_6344 & _T_7830; // @[LoadQueue.scala 131:72:@8813.4]
  assign _T_7833 = offsetQ_0 < 4'hd; // @[LoadQueue.scala 132:33:@8814.4]
  assign _T_7836 = _T_7833 & _T_6353; // @[LoadQueue.scala 132:41:@8816.4]
  assign _T_7838 = _T_7836 == 1'h0; // @[LoadQueue.scala 132:9:@8817.4]
  assign storesToCheck_0_13 = _T_2236 ? _T_7831 : _T_7838; // @[LoadQueue.scala 131:10:@8818.4]
  assign _T_7844 = 4'he <= offsetQ_0; // @[LoadQueue.scala 131:81:@8821.4]
  assign _T_7845 = _T_6361 & _T_7844; // @[LoadQueue.scala 131:72:@8822.4]
  assign _T_7847 = offsetQ_0 < 4'he; // @[LoadQueue.scala 132:33:@8823.4]
  assign _T_7850 = _T_7847 & _T_6370; // @[LoadQueue.scala 132:41:@8825.4]
  assign _T_7852 = _T_7850 == 1'h0; // @[LoadQueue.scala 132:9:@8826.4]
  assign storesToCheck_0_14 = _T_2236 ? _T_7845 : _T_7852; // @[LoadQueue.scala 131:10:@8827.4]
  assign _T_7858 = 4'hf <= offsetQ_0; // @[LoadQueue.scala 131:81:@8830.4]
  assign storesToCheck_0_15 = _T_2236 ? _T_7858 : 1'h1; // @[LoadQueue.scala 131:10:@8836.4]
  assign storesToCheck_1_0 = _T_2266 ? _T_6123 : 1'h1; // @[LoadQueue.scala 131:10:@8878.4]
  assign _T_7908 = 4'h1 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8881.4]
  assign _T_7909 = _T_6140 & _T_7908; // @[LoadQueue.scala 131:72:@8882.4]
  assign _T_7911 = offsetQ_1 < 4'h1; // @[LoadQueue.scala 132:33:@8883.4]
  assign _T_7914 = _T_7911 & _T_6149; // @[LoadQueue.scala 132:41:@8885.4]
  assign _T_7916 = _T_7914 == 1'h0; // @[LoadQueue.scala 132:9:@8886.4]
  assign storesToCheck_1_1 = _T_2266 ? _T_7909 : _T_7916; // @[LoadQueue.scala 131:10:@8887.4]
  assign _T_7922 = 4'h2 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8890.4]
  assign _T_7923 = _T_6157 & _T_7922; // @[LoadQueue.scala 131:72:@8891.4]
  assign _T_7925 = offsetQ_1 < 4'h2; // @[LoadQueue.scala 132:33:@8892.4]
  assign _T_7928 = _T_7925 & _T_6166; // @[LoadQueue.scala 132:41:@8894.4]
  assign _T_7930 = _T_7928 == 1'h0; // @[LoadQueue.scala 132:9:@8895.4]
  assign storesToCheck_1_2 = _T_2266 ? _T_7923 : _T_7930; // @[LoadQueue.scala 131:10:@8896.4]
  assign _T_7936 = 4'h3 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8899.4]
  assign _T_7937 = _T_6174 & _T_7936; // @[LoadQueue.scala 131:72:@8900.4]
  assign _T_7939 = offsetQ_1 < 4'h3; // @[LoadQueue.scala 132:33:@8901.4]
  assign _T_7942 = _T_7939 & _T_6183; // @[LoadQueue.scala 132:41:@8903.4]
  assign _T_7944 = _T_7942 == 1'h0; // @[LoadQueue.scala 132:9:@8904.4]
  assign storesToCheck_1_3 = _T_2266 ? _T_7937 : _T_7944; // @[LoadQueue.scala 131:10:@8905.4]
  assign _T_7950 = 4'h4 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8908.4]
  assign _T_7951 = _T_6191 & _T_7950; // @[LoadQueue.scala 131:72:@8909.4]
  assign _T_7953 = offsetQ_1 < 4'h4; // @[LoadQueue.scala 132:33:@8910.4]
  assign _T_7956 = _T_7953 & _T_6200; // @[LoadQueue.scala 132:41:@8912.4]
  assign _T_7958 = _T_7956 == 1'h0; // @[LoadQueue.scala 132:9:@8913.4]
  assign storesToCheck_1_4 = _T_2266 ? _T_7951 : _T_7958; // @[LoadQueue.scala 131:10:@8914.4]
  assign _T_7964 = 4'h5 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8917.4]
  assign _T_7965 = _T_6208 & _T_7964; // @[LoadQueue.scala 131:72:@8918.4]
  assign _T_7967 = offsetQ_1 < 4'h5; // @[LoadQueue.scala 132:33:@8919.4]
  assign _T_7970 = _T_7967 & _T_6217; // @[LoadQueue.scala 132:41:@8921.4]
  assign _T_7972 = _T_7970 == 1'h0; // @[LoadQueue.scala 132:9:@8922.4]
  assign storesToCheck_1_5 = _T_2266 ? _T_7965 : _T_7972; // @[LoadQueue.scala 131:10:@8923.4]
  assign _T_7978 = 4'h6 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8926.4]
  assign _T_7979 = _T_6225 & _T_7978; // @[LoadQueue.scala 131:72:@8927.4]
  assign _T_7981 = offsetQ_1 < 4'h6; // @[LoadQueue.scala 132:33:@8928.4]
  assign _T_7984 = _T_7981 & _T_6234; // @[LoadQueue.scala 132:41:@8930.4]
  assign _T_7986 = _T_7984 == 1'h0; // @[LoadQueue.scala 132:9:@8931.4]
  assign storesToCheck_1_6 = _T_2266 ? _T_7979 : _T_7986; // @[LoadQueue.scala 131:10:@8932.4]
  assign _T_7992 = 4'h7 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8935.4]
  assign _T_7993 = _T_6242 & _T_7992; // @[LoadQueue.scala 131:72:@8936.4]
  assign _T_7995 = offsetQ_1 < 4'h7; // @[LoadQueue.scala 132:33:@8937.4]
  assign _T_7998 = _T_7995 & _T_6251; // @[LoadQueue.scala 132:41:@8939.4]
  assign _T_8000 = _T_7998 == 1'h0; // @[LoadQueue.scala 132:9:@8940.4]
  assign storesToCheck_1_7 = _T_2266 ? _T_7993 : _T_8000; // @[LoadQueue.scala 131:10:@8941.4]
  assign _T_8006 = 4'h8 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8944.4]
  assign _T_8007 = _T_6259 & _T_8006; // @[LoadQueue.scala 131:72:@8945.4]
  assign _T_8009 = offsetQ_1 < 4'h8; // @[LoadQueue.scala 132:33:@8946.4]
  assign _T_8012 = _T_8009 & _T_6268; // @[LoadQueue.scala 132:41:@8948.4]
  assign _T_8014 = _T_8012 == 1'h0; // @[LoadQueue.scala 132:9:@8949.4]
  assign storesToCheck_1_8 = _T_2266 ? _T_8007 : _T_8014; // @[LoadQueue.scala 131:10:@8950.4]
  assign _T_8020 = 4'h9 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8953.4]
  assign _T_8021 = _T_6276 & _T_8020; // @[LoadQueue.scala 131:72:@8954.4]
  assign _T_8023 = offsetQ_1 < 4'h9; // @[LoadQueue.scala 132:33:@8955.4]
  assign _T_8026 = _T_8023 & _T_6285; // @[LoadQueue.scala 132:41:@8957.4]
  assign _T_8028 = _T_8026 == 1'h0; // @[LoadQueue.scala 132:9:@8958.4]
  assign storesToCheck_1_9 = _T_2266 ? _T_8021 : _T_8028; // @[LoadQueue.scala 131:10:@8959.4]
  assign _T_8034 = 4'ha <= offsetQ_1; // @[LoadQueue.scala 131:81:@8962.4]
  assign _T_8035 = _T_6293 & _T_8034; // @[LoadQueue.scala 131:72:@8963.4]
  assign _T_8037 = offsetQ_1 < 4'ha; // @[LoadQueue.scala 132:33:@8964.4]
  assign _T_8040 = _T_8037 & _T_6302; // @[LoadQueue.scala 132:41:@8966.4]
  assign _T_8042 = _T_8040 == 1'h0; // @[LoadQueue.scala 132:9:@8967.4]
  assign storesToCheck_1_10 = _T_2266 ? _T_8035 : _T_8042; // @[LoadQueue.scala 131:10:@8968.4]
  assign _T_8048 = 4'hb <= offsetQ_1; // @[LoadQueue.scala 131:81:@8971.4]
  assign _T_8049 = _T_6310 & _T_8048; // @[LoadQueue.scala 131:72:@8972.4]
  assign _T_8051 = offsetQ_1 < 4'hb; // @[LoadQueue.scala 132:33:@8973.4]
  assign _T_8054 = _T_8051 & _T_6319; // @[LoadQueue.scala 132:41:@8975.4]
  assign _T_8056 = _T_8054 == 1'h0; // @[LoadQueue.scala 132:9:@8976.4]
  assign storesToCheck_1_11 = _T_2266 ? _T_8049 : _T_8056; // @[LoadQueue.scala 131:10:@8977.4]
  assign _T_8062 = 4'hc <= offsetQ_1; // @[LoadQueue.scala 131:81:@8980.4]
  assign _T_8063 = _T_6327 & _T_8062; // @[LoadQueue.scala 131:72:@8981.4]
  assign _T_8065 = offsetQ_1 < 4'hc; // @[LoadQueue.scala 132:33:@8982.4]
  assign _T_8068 = _T_8065 & _T_6336; // @[LoadQueue.scala 132:41:@8984.4]
  assign _T_8070 = _T_8068 == 1'h0; // @[LoadQueue.scala 132:9:@8985.4]
  assign storesToCheck_1_12 = _T_2266 ? _T_8063 : _T_8070; // @[LoadQueue.scala 131:10:@8986.4]
  assign _T_8076 = 4'hd <= offsetQ_1; // @[LoadQueue.scala 131:81:@8989.4]
  assign _T_8077 = _T_6344 & _T_8076; // @[LoadQueue.scala 131:72:@8990.4]
  assign _T_8079 = offsetQ_1 < 4'hd; // @[LoadQueue.scala 132:33:@8991.4]
  assign _T_8082 = _T_8079 & _T_6353; // @[LoadQueue.scala 132:41:@8993.4]
  assign _T_8084 = _T_8082 == 1'h0; // @[LoadQueue.scala 132:9:@8994.4]
  assign storesToCheck_1_13 = _T_2266 ? _T_8077 : _T_8084; // @[LoadQueue.scala 131:10:@8995.4]
  assign _T_8090 = 4'he <= offsetQ_1; // @[LoadQueue.scala 131:81:@8998.4]
  assign _T_8091 = _T_6361 & _T_8090; // @[LoadQueue.scala 131:72:@8999.4]
  assign _T_8093 = offsetQ_1 < 4'he; // @[LoadQueue.scala 132:33:@9000.4]
  assign _T_8096 = _T_8093 & _T_6370; // @[LoadQueue.scala 132:41:@9002.4]
  assign _T_8098 = _T_8096 == 1'h0; // @[LoadQueue.scala 132:9:@9003.4]
  assign storesToCheck_1_14 = _T_2266 ? _T_8091 : _T_8098; // @[LoadQueue.scala 131:10:@9004.4]
  assign _T_8104 = 4'hf <= offsetQ_1; // @[LoadQueue.scala 131:81:@9007.4]
  assign storesToCheck_1_15 = _T_2266 ? _T_8104 : 1'h1; // @[LoadQueue.scala 131:10:@9013.4]
  assign storesToCheck_2_0 = _T_2296 ? _T_6123 : 1'h1; // @[LoadQueue.scala 131:10:@9055.4]
  assign _T_8154 = 4'h1 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9058.4]
  assign _T_8155 = _T_6140 & _T_8154; // @[LoadQueue.scala 131:72:@9059.4]
  assign _T_8157 = offsetQ_2 < 4'h1; // @[LoadQueue.scala 132:33:@9060.4]
  assign _T_8160 = _T_8157 & _T_6149; // @[LoadQueue.scala 132:41:@9062.4]
  assign _T_8162 = _T_8160 == 1'h0; // @[LoadQueue.scala 132:9:@9063.4]
  assign storesToCheck_2_1 = _T_2296 ? _T_8155 : _T_8162; // @[LoadQueue.scala 131:10:@9064.4]
  assign _T_8168 = 4'h2 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9067.4]
  assign _T_8169 = _T_6157 & _T_8168; // @[LoadQueue.scala 131:72:@9068.4]
  assign _T_8171 = offsetQ_2 < 4'h2; // @[LoadQueue.scala 132:33:@9069.4]
  assign _T_8174 = _T_8171 & _T_6166; // @[LoadQueue.scala 132:41:@9071.4]
  assign _T_8176 = _T_8174 == 1'h0; // @[LoadQueue.scala 132:9:@9072.4]
  assign storesToCheck_2_2 = _T_2296 ? _T_8169 : _T_8176; // @[LoadQueue.scala 131:10:@9073.4]
  assign _T_8182 = 4'h3 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9076.4]
  assign _T_8183 = _T_6174 & _T_8182; // @[LoadQueue.scala 131:72:@9077.4]
  assign _T_8185 = offsetQ_2 < 4'h3; // @[LoadQueue.scala 132:33:@9078.4]
  assign _T_8188 = _T_8185 & _T_6183; // @[LoadQueue.scala 132:41:@9080.4]
  assign _T_8190 = _T_8188 == 1'h0; // @[LoadQueue.scala 132:9:@9081.4]
  assign storesToCheck_2_3 = _T_2296 ? _T_8183 : _T_8190; // @[LoadQueue.scala 131:10:@9082.4]
  assign _T_8196 = 4'h4 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9085.4]
  assign _T_8197 = _T_6191 & _T_8196; // @[LoadQueue.scala 131:72:@9086.4]
  assign _T_8199 = offsetQ_2 < 4'h4; // @[LoadQueue.scala 132:33:@9087.4]
  assign _T_8202 = _T_8199 & _T_6200; // @[LoadQueue.scala 132:41:@9089.4]
  assign _T_8204 = _T_8202 == 1'h0; // @[LoadQueue.scala 132:9:@9090.4]
  assign storesToCheck_2_4 = _T_2296 ? _T_8197 : _T_8204; // @[LoadQueue.scala 131:10:@9091.4]
  assign _T_8210 = 4'h5 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9094.4]
  assign _T_8211 = _T_6208 & _T_8210; // @[LoadQueue.scala 131:72:@9095.4]
  assign _T_8213 = offsetQ_2 < 4'h5; // @[LoadQueue.scala 132:33:@9096.4]
  assign _T_8216 = _T_8213 & _T_6217; // @[LoadQueue.scala 132:41:@9098.4]
  assign _T_8218 = _T_8216 == 1'h0; // @[LoadQueue.scala 132:9:@9099.4]
  assign storesToCheck_2_5 = _T_2296 ? _T_8211 : _T_8218; // @[LoadQueue.scala 131:10:@9100.4]
  assign _T_8224 = 4'h6 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9103.4]
  assign _T_8225 = _T_6225 & _T_8224; // @[LoadQueue.scala 131:72:@9104.4]
  assign _T_8227 = offsetQ_2 < 4'h6; // @[LoadQueue.scala 132:33:@9105.4]
  assign _T_8230 = _T_8227 & _T_6234; // @[LoadQueue.scala 132:41:@9107.4]
  assign _T_8232 = _T_8230 == 1'h0; // @[LoadQueue.scala 132:9:@9108.4]
  assign storesToCheck_2_6 = _T_2296 ? _T_8225 : _T_8232; // @[LoadQueue.scala 131:10:@9109.4]
  assign _T_8238 = 4'h7 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9112.4]
  assign _T_8239 = _T_6242 & _T_8238; // @[LoadQueue.scala 131:72:@9113.4]
  assign _T_8241 = offsetQ_2 < 4'h7; // @[LoadQueue.scala 132:33:@9114.4]
  assign _T_8244 = _T_8241 & _T_6251; // @[LoadQueue.scala 132:41:@9116.4]
  assign _T_8246 = _T_8244 == 1'h0; // @[LoadQueue.scala 132:9:@9117.4]
  assign storesToCheck_2_7 = _T_2296 ? _T_8239 : _T_8246; // @[LoadQueue.scala 131:10:@9118.4]
  assign _T_8252 = 4'h8 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9121.4]
  assign _T_8253 = _T_6259 & _T_8252; // @[LoadQueue.scala 131:72:@9122.4]
  assign _T_8255 = offsetQ_2 < 4'h8; // @[LoadQueue.scala 132:33:@9123.4]
  assign _T_8258 = _T_8255 & _T_6268; // @[LoadQueue.scala 132:41:@9125.4]
  assign _T_8260 = _T_8258 == 1'h0; // @[LoadQueue.scala 132:9:@9126.4]
  assign storesToCheck_2_8 = _T_2296 ? _T_8253 : _T_8260; // @[LoadQueue.scala 131:10:@9127.4]
  assign _T_8266 = 4'h9 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9130.4]
  assign _T_8267 = _T_6276 & _T_8266; // @[LoadQueue.scala 131:72:@9131.4]
  assign _T_8269 = offsetQ_2 < 4'h9; // @[LoadQueue.scala 132:33:@9132.4]
  assign _T_8272 = _T_8269 & _T_6285; // @[LoadQueue.scala 132:41:@9134.4]
  assign _T_8274 = _T_8272 == 1'h0; // @[LoadQueue.scala 132:9:@9135.4]
  assign storesToCheck_2_9 = _T_2296 ? _T_8267 : _T_8274; // @[LoadQueue.scala 131:10:@9136.4]
  assign _T_8280 = 4'ha <= offsetQ_2; // @[LoadQueue.scala 131:81:@9139.4]
  assign _T_8281 = _T_6293 & _T_8280; // @[LoadQueue.scala 131:72:@9140.4]
  assign _T_8283 = offsetQ_2 < 4'ha; // @[LoadQueue.scala 132:33:@9141.4]
  assign _T_8286 = _T_8283 & _T_6302; // @[LoadQueue.scala 132:41:@9143.4]
  assign _T_8288 = _T_8286 == 1'h0; // @[LoadQueue.scala 132:9:@9144.4]
  assign storesToCheck_2_10 = _T_2296 ? _T_8281 : _T_8288; // @[LoadQueue.scala 131:10:@9145.4]
  assign _T_8294 = 4'hb <= offsetQ_2; // @[LoadQueue.scala 131:81:@9148.4]
  assign _T_8295 = _T_6310 & _T_8294; // @[LoadQueue.scala 131:72:@9149.4]
  assign _T_8297 = offsetQ_2 < 4'hb; // @[LoadQueue.scala 132:33:@9150.4]
  assign _T_8300 = _T_8297 & _T_6319; // @[LoadQueue.scala 132:41:@9152.4]
  assign _T_8302 = _T_8300 == 1'h0; // @[LoadQueue.scala 132:9:@9153.4]
  assign storesToCheck_2_11 = _T_2296 ? _T_8295 : _T_8302; // @[LoadQueue.scala 131:10:@9154.4]
  assign _T_8308 = 4'hc <= offsetQ_2; // @[LoadQueue.scala 131:81:@9157.4]
  assign _T_8309 = _T_6327 & _T_8308; // @[LoadQueue.scala 131:72:@9158.4]
  assign _T_8311 = offsetQ_2 < 4'hc; // @[LoadQueue.scala 132:33:@9159.4]
  assign _T_8314 = _T_8311 & _T_6336; // @[LoadQueue.scala 132:41:@9161.4]
  assign _T_8316 = _T_8314 == 1'h0; // @[LoadQueue.scala 132:9:@9162.4]
  assign storesToCheck_2_12 = _T_2296 ? _T_8309 : _T_8316; // @[LoadQueue.scala 131:10:@9163.4]
  assign _T_8322 = 4'hd <= offsetQ_2; // @[LoadQueue.scala 131:81:@9166.4]
  assign _T_8323 = _T_6344 & _T_8322; // @[LoadQueue.scala 131:72:@9167.4]
  assign _T_8325 = offsetQ_2 < 4'hd; // @[LoadQueue.scala 132:33:@9168.4]
  assign _T_8328 = _T_8325 & _T_6353; // @[LoadQueue.scala 132:41:@9170.4]
  assign _T_8330 = _T_8328 == 1'h0; // @[LoadQueue.scala 132:9:@9171.4]
  assign storesToCheck_2_13 = _T_2296 ? _T_8323 : _T_8330; // @[LoadQueue.scala 131:10:@9172.4]
  assign _T_8336 = 4'he <= offsetQ_2; // @[LoadQueue.scala 131:81:@9175.4]
  assign _T_8337 = _T_6361 & _T_8336; // @[LoadQueue.scala 131:72:@9176.4]
  assign _T_8339 = offsetQ_2 < 4'he; // @[LoadQueue.scala 132:33:@9177.4]
  assign _T_8342 = _T_8339 & _T_6370; // @[LoadQueue.scala 132:41:@9179.4]
  assign _T_8344 = _T_8342 == 1'h0; // @[LoadQueue.scala 132:9:@9180.4]
  assign storesToCheck_2_14 = _T_2296 ? _T_8337 : _T_8344; // @[LoadQueue.scala 131:10:@9181.4]
  assign _T_8350 = 4'hf <= offsetQ_2; // @[LoadQueue.scala 131:81:@9184.4]
  assign storesToCheck_2_15 = _T_2296 ? _T_8350 : 1'h1; // @[LoadQueue.scala 131:10:@9190.4]
  assign storesToCheck_3_0 = _T_2326 ? _T_6123 : 1'h1; // @[LoadQueue.scala 131:10:@9232.4]
  assign _T_8400 = 4'h1 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9235.4]
  assign _T_8401 = _T_6140 & _T_8400; // @[LoadQueue.scala 131:72:@9236.4]
  assign _T_8403 = offsetQ_3 < 4'h1; // @[LoadQueue.scala 132:33:@9237.4]
  assign _T_8406 = _T_8403 & _T_6149; // @[LoadQueue.scala 132:41:@9239.4]
  assign _T_8408 = _T_8406 == 1'h0; // @[LoadQueue.scala 132:9:@9240.4]
  assign storesToCheck_3_1 = _T_2326 ? _T_8401 : _T_8408; // @[LoadQueue.scala 131:10:@9241.4]
  assign _T_8414 = 4'h2 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9244.4]
  assign _T_8415 = _T_6157 & _T_8414; // @[LoadQueue.scala 131:72:@9245.4]
  assign _T_8417 = offsetQ_3 < 4'h2; // @[LoadQueue.scala 132:33:@9246.4]
  assign _T_8420 = _T_8417 & _T_6166; // @[LoadQueue.scala 132:41:@9248.4]
  assign _T_8422 = _T_8420 == 1'h0; // @[LoadQueue.scala 132:9:@9249.4]
  assign storesToCheck_3_2 = _T_2326 ? _T_8415 : _T_8422; // @[LoadQueue.scala 131:10:@9250.4]
  assign _T_8428 = 4'h3 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9253.4]
  assign _T_8429 = _T_6174 & _T_8428; // @[LoadQueue.scala 131:72:@9254.4]
  assign _T_8431 = offsetQ_3 < 4'h3; // @[LoadQueue.scala 132:33:@9255.4]
  assign _T_8434 = _T_8431 & _T_6183; // @[LoadQueue.scala 132:41:@9257.4]
  assign _T_8436 = _T_8434 == 1'h0; // @[LoadQueue.scala 132:9:@9258.4]
  assign storesToCheck_3_3 = _T_2326 ? _T_8429 : _T_8436; // @[LoadQueue.scala 131:10:@9259.4]
  assign _T_8442 = 4'h4 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9262.4]
  assign _T_8443 = _T_6191 & _T_8442; // @[LoadQueue.scala 131:72:@9263.4]
  assign _T_8445 = offsetQ_3 < 4'h4; // @[LoadQueue.scala 132:33:@9264.4]
  assign _T_8448 = _T_8445 & _T_6200; // @[LoadQueue.scala 132:41:@9266.4]
  assign _T_8450 = _T_8448 == 1'h0; // @[LoadQueue.scala 132:9:@9267.4]
  assign storesToCheck_3_4 = _T_2326 ? _T_8443 : _T_8450; // @[LoadQueue.scala 131:10:@9268.4]
  assign _T_8456 = 4'h5 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9271.4]
  assign _T_8457 = _T_6208 & _T_8456; // @[LoadQueue.scala 131:72:@9272.4]
  assign _T_8459 = offsetQ_3 < 4'h5; // @[LoadQueue.scala 132:33:@9273.4]
  assign _T_8462 = _T_8459 & _T_6217; // @[LoadQueue.scala 132:41:@9275.4]
  assign _T_8464 = _T_8462 == 1'h0; // @[LoadQueue.scala 132:9:@9276.4]
  assign storesToCheck_3_5 = _T_2326 ? _T_8457 : _T_8464; // @[LoadQueue.scala 131:10:@9277.4]
  assign _T_8470 = 4'h6 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9280.4]
  assign _T_8471 = _T_6225 & _T_8470; // @[LoadQueue.scala 131:72:@9281.4]
  assign _T_8473 = offsetQ_3 < 4'h6; // @[LoadQueue.scala 132:33:@9282.4]
  assign _T_8476 = _T_8473 & _T_6234; // @[LoadQueue.scala 132:41:@9284.4]
  assign _T_8478 = _T_8476 == 1'h0; // @[LoadQueue.scala 132:9:@9285.4]
  assign storesToCheck_3_6 = _T_2326 ? _T_8471 : _T_8478; // @[LoadQueue.scala 131:10:@9286.4]
  assign _T_8484 = 4'h7 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9289.4]
  assign _T_8485 = _T_6242 & _T_8484; // @[LoadQueue.scala 131:72:@9290.4]
  assign _T_8487 = offsetQ_3 < 4'h7; // @[LoadQueue.scala 132:33:@9291.4]
  assign _T_8490 = _T_8487 & _T_6251; // @[LoadQueue.scala 132:41:@9293.4]
  assign _T_8492 = _T_8490 == 1'h0; // @[LoadQueue.scala 132:9:@9294.4]
  assign storesToCheck_3_7 = _T_2326 ? _T_8485 : _T_8492; // @[LoadQueue.scala 131:10:@9295.4]
  assign _T_8498 = 4'h8 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9298.4]
  assign _T_8499 = _T_6259 & _T_8498; // @[LoadQueue.scala 131:72:@9299.4]
  assign _T_8501 = offsetQ_3 < 4'h8; // @[LoadQueue.scala 132:33:@9300.4]
  assign _T_8504 = _T_8501 & _T_6268; // @[LoadQueue.scala 132:41:@9302.4]
  assign _T_8506 = _T_8504 == 1'h0; // @[LoadQueue.scala 132:9:@9303.4]
  assign storesToCheck_3_8 = _T_2326 ? _T_8499 : _T_8506; // @[LoadQueue.scala 131:10:@9304.4]
  assign _T_8512 = 4'h9 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9307.4]
  assign _T_8513 = _T_6276 & _T_8512; // @[LoadQueue.scala 131:72:@9308.4]
  assign _T_8515 = offsetQ_3 < 4'h9; // @[LoadQueue.scala 132:33:@9309.4]
  assign _T_8518 = _T_8515 & _T_6285; // @[LoadQueue.scala 132:41:@9311.4]
  assign _T_8520 = _T_8518 == 1'h0; // @[LoadQueue.scala 132:9:@9312.4]
  assign storesToCheck_3_9 = _T_2326 ? _T_8513 : _T_8520; // @[LoadQueue.scala 131:10:@9313.4]
  assign _T_8526 = 4'ha <= offsetQ_3; // @[LoadQueue.scala 131:81:@9316.4]
  assign _T_8527 = _T_6293 & _T_8526; // @[LoadQueue.scala 131:72:@9317.4]
  assign _T_8529 = offsetQ_3 < 4'ha; // @[LoadQueue.scala 132:33:@9318.4]
  assign _T_8532 = _T_8529 & _T_6302; // @[LoadQueue.scala 132:41:@9320.4]
  assign _T_8534 = _T_8532 == 1'h0; // @[LoadQueue.scala 132:9:@9321.4]
  assign storesToCheck_3_10 = _T_2326 ? _T_8527 : _T_8534; // @[LoadQueue.scala 131:10:@9322.4]
  assign _T_8540 = 4'hb <= offsetQ_3; // @[LoadQueue.scala 131:81:@9325.4]
  assign _T_8541 = _T_6310 & _T_8540; // @[LoadQueue.scala 131:72:@9326.4]
  assign _T_8543 = offsetQ_3 < 4'hb; // @[LoadQueue.scala 132:33:@9327.4]
  assign _T_8546 = _T_8543 & _T_6319; // @[LoadQueue.scala 132:41:@9329.4]
  assign _T_8548 = _T_8546 == 1'h0; // @[LoadQueue.scala 132:9:@9330.4]
  assign storesToCheck_3_11 = _T_2326 ? _T_8541 : _T_8548; // @[LoadQueue.scala 131:10:@9331.4]
  assign _T_8554 = 4'hc <= offsetQ_3; // @[LoadQueue.scala 131:81:@9334.4]
  assign _T_8555 = _T_6327 & _T_8554; // @[LoadQueue.scala 131:72:@9335.4]
  assign _T_8557 = offsetQ_3 < 4'hc; // @[LoadQueue.scala 132:33:@9336.4]
  assign _T_8560 = _T_8557 & _T_6336; // @[LoadQueue.scala 132:41:@9338.4]
  assign _T_8562 = _T_8560 == 1'h0; // @[LoadQueue.scala 132:9:@9339.4]
  assign storesToCheck_3_12 = _T_2326 ? _T_8555 : _T_8562; // @[LoadQueue.scala 131:10:@9340.4]
  assign _T_8568 = 4'hd <= offsetQ_3; // @[LoadQueue.scala 131:81:@9343.4]
  assign _T_8569 = _T_6344 & _T_8568; // @[LoadQueue.scala 131:72:@9344.4]
  assign _T_8571 = offsetQ_3 < 4'hd; // @[LoadQueue.scala 132:33:@9345.4]
  assign _T_8574 = _T_8571 & _T_6353; // @[LoadQueue.scala 132:41:@9347.4]
  assign _T_8576 = _T_8574 == 1'h0; // @[LoadQueue.scala 132:9:@9348.4]
  assign storesToCheck_3_13 = _T_2326 ? _T_8569 : _T_8576; // @[LoadQueue.scala 131:10:@9349.4]
  assign _T_8582 = 4'he <= offsetQ_3; // @[LoadQueue.scala 131:81:@9352.4]
  assign _T_8583 = _T_6361 & _T_8582; // @[LoadQueue.scala 131:72:@9353.4]
  assign _T_8585 = offsetQ_3 < 4'he; // @[LoadQueue.scala 132:33:@9354.4]
  assign _T_8588 = _T_8585 & _T_6370; // @[LoadQueue.scala 132:41:@9356.4]
  assign _T_8590 = _T_8588 == 1'h0; // @[LoadQueue.scala 132:9:@9357.4]
  assign storesToCheck_3_14 = _T_2326 ? _T_8583 : _T_8590; // @[LoadQueue.scala 131:10:@9358.4]
  assign _T_8596 = 4'hf <= offsetQ_3; // @[LoadQueue.scala 131:81:@9361.4]
  assign storesToCheck_3_15 = _T_2326 ? _T_8596 : 1'h1; // @[LoadQueue.scala 131:10:@9367.4]
  assign storesToCheck_4_0 = _T_2356 ? _T_6123 : 1'h1; // @[LoadQueue.scala 131:10:@9409.4]
  assign _T_8646 = 4'h1 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9412.4]
  assign _T_8647 = _T_6140 & _T_8646; // @[LoadQueue.scala 131:72:@9413.4]
  assign _T_8649 = offsetQ_4 < 4'h1; // @[LoadQueue.scala 132:33:@9414.4]
  assign _T_8652 = _T_8649 & _T_6149; // @[LoadQueue.scala 132:41:@9416.4]
  assign _T_8654 = _T_8652 == 1'h0; // @[LoadQueue.scala 132:9:@9417.4]
  assign storesToCheck_4_1 = _T_2356 ? _T_8647 : _T_8654; // @[LoadQueue.scala 131:10:@9418.4]
  assign _T_8660 = 4'h2 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9421.4]
  assign _T_8661 = _T_6157 & _T_8660; // @[LoadQueue.scala 131:72:@9422.4]
  assign _T_8663 = offsetQ_4 < 4'h2; // @[LoadQueue.scala 132:33:@9423.4]
  assign _T_8666 = _T_8663 & _T_6166; // @[LoadQueue.scala 132:41:@9425.4]
  assign _T_8668 = _T_8666 == 1'h0; // @[LoadQueue.scala 132:9:@9426.4]
  assign storesToCheck_4_2 = _T_2356 ? _T_8661 : _T_8668; // @[LoadQueue.scala 131:10:@9427.4]
  assign _T_8674 = 4'h3 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9430.4]
  assign _T_8675 = _T_6174 & _T_8674; // @[LoadQueue.scala 131:72:@9431.4]
  assign _T_8677 = offsetQ_4 < 4'h3; // @[LoadQueue.scala 132:33:@9432.4]
  assign _T_8680 = _T_8677 & _T_6183; // @[LoadQueue.scala 132:41:@9434.4]
  assign _T_8682 = _T_8680 == 1'h0; // @[LoadQueue.scala 132:9:@9435.4]
  assign storesToCheck_4_3 = _T_2356 ? _T_8675 : _T_8682; // @[LoadQueue.scala 131:10:@9436.4]
  assign _T_8688 = 4'h4 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9439.4]
  assign _T_8689 = _T_6191 & _T_8688; // @[LoadQueue.scala 131:72:@9440.4]
  assign _T_8691 = offsetQ_4 < 4'h4; // @[LoadQueue.scala 132:33:@9441.4]
  assign _T_8694 = _T_8691 & _T_6200; // @[LoadQueue.scala 132:41:@9443.4]
  assign _T_8696 = _T_8694 == 1'h0; // @[LoadQueue.scala 132:9:@9444.4]
  assign storesToCheck_4_4 = _T_2356 ? _T_8689 : _T_8696; // @[LoadQueue.scala 131:10:@9445.4]
  assign _T_8702 = 4'h5 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9448.4]
  assign _T_8703 = _T_6208 & _T_8702; // @[LoadQueue.scala 131:72:@9449.4]
  assign _T_8705 = offsetQ_4 < 4'h5; // @[LoadQueue.scala 132:33:@9450.4]
  assign _T_8708 = _T_8705 & _T_6217; // @[LoadQueue.scala 132:41:@9452.4]
  assign _T_8710 = _T_8708 == 1'h0; // @[LoadQueue.scala 132:9:@9453.4]
  assign storesToCheck_4_5 = _T_2356 ? _T_8703 : _T_8710; // @[LoadQueue.scala 131:10:@9454.4]
  assign _T_8716 = 4'h6 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9457.4]
  assign _T_8717 = _T_6225 & _T_8716; // @[LoadQueue.scala 131:72:@9458.4]
  assign _T_8719 = offsetQ_4 < 4'h6; // @[LoadQueue.scala 132:33:@9459.4]
  assign _T_8722 = _T_8719 & _T_6234; // @[LoadQueue.scala 132:41:@9461.4]
  assign _T_8724 = _T_8722 == 1'h0; // @[LoadQueue.scala 132:9:@9462.4]
  assign storesToCheck_4_6 = _T_2356 ? _T_8717 : _T_8724; // @[LoadQueue.scala 131:10:@9463.4]
  assign _T_8730 = 4'h7 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9466.4]
  assign _T_8731 = _T_6242 & _T_8730; // @[LoadQueue.scala 131:72:@9467.4]
  assign _T_8733 = offsetQ_4 < 4'h7; // @[LoadQueue.scala 132:33:@9468.4]
  assign _T_8736 = _T_8733 & _T_6251; // @[LoadQueue.scala 132:41:@9470.4]
  assign _T_8738 = _T_8736 == 1'h0; // @[LoadQueue.scala 132:9:@9471.4]
  assign storesToCheck_4_7 = _T_2356 ? _T_8731 : _T_8738; // @[LoadQueue.scala 131:10:@9472.4]
  assign _T_8744 = 4'h8 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9475.4]
  assign _T_8745 = _T_6259 & _T_8744; // @[LoadQueue.scala 131:72:@9476.4]
  assign _T_8747 = offsetQ_4 < 4'h8; // @[LoadQueue.scala 132:33:@9477.4]
  assign _T_8750 = _T_8747 & _T_6268; // @[LoadQueue.scala 132:41:@9479.4]
  assign _T_8752 = _T_8750 == 1'h0; // @[LoadQueue.scala 132:9:@9480.4]
  assign storesToCheck_4_8 = _T_2356 ? _T_8745 : _T_8752; // @[LoadQueue.scala 131:10:@9481.4]
  assign _T_8758 = 4'h9 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9484.4]
  assign _T_8759 = _T_6276 & _T_8758; // @[LoadQueue.scala 131:72:@9485.4]
  assign _T_8761 = offsetQ_4 < 4'h9; // @[LoadQueue.scala 132:33:@9486.4]
  assign _T_8764 = _T_8761 & _T_6285; // @[LoadQueue.scala 132:41:@9488.4]
  assign _T_8766 = _T_8764 == 1'h0; // @[LoadQueue.scala 132:9:@9489.4]
  assign storesToCheck_4_9 = _T_2356 ? _T_8759 : _T_8766; // @[LoadQueue.scala 131:10:@9490.4]
  assign _T_8772 = 4'ha <= offsetQ_4; // @[LoadQueue.scala 131:81:@9493.4]
  assign _T_8773 = _T_6293 & _T_8772; // @[LoadQueue.scala 131:72:@9494.4]
  assign _T_8775 = offsetQ_4 < 4'ha; // @[LoadQueue.scala 132:33:@9495.4]
  assign _T_8778 = _T_8775 & _T_6302; // @[LoadQueue.scala 132:41:@9497.4]
  assign _T_8780 = _T_8778 == 1'h0; // @[LoadQueue.scala 132:9:@9498.4]
  assign storesToCheck_4_10 = _T_2356 ? _T_8773 : _T_8780; // @[LoadQueue.scala 131:10:@9499.4]
  assign _T_8786 = 4'hb <= offsetQ_4; // @[LoadQueue.scala 131:81:@9502.4]
  assign _T_8787 = _T_6310 & _T_8786; // @[LoadQueue.scala 131:72:@9503.4]
  assign _T_8789 = offsetQ_4 < 4'hb; // @[LoadQueue.scala 132:33:@9504.4]
  assign _T_8792 = _T_8789 & _T_6319; // @[LoadQueue.scala 132:41:@9506.4]
  assign _T_8794 = _T_8792 == 1'h0; // @[LoadQueue.scala 132:9:@9507.4]
  assign storesToCheck_4_11 = _T_2356 ? _T_8787 : _T_8794; // @[LoadQueue.scala 131:10:@9508.4]
  assign _T_8800 = 4'hc <= offsetQ_4; // @[LoadQueue.scala 131:81:@9511.4]
  assign _T_8801 = _T_6327 & _T_8800; // @[LoadQueue.scala 131:72:@9512.4]
  assign _T_8803 = offsetQ_4 < 4'hc; // @[LoadQueue.scala 132:33:@9513.4]
  assign _T_8806 = _T_8803 & _T_6336; // @[LoadQueue.scala 132:41:@9515.4]
  assign _T_8808 = _T_8806 == 1'h0; // @[LoadQueue.scala 132:9:@9516.4]
  assign storesToCheck_4_12 = _T_2356 ? _T_8801 : _T_8808; // @[LoadQueue.scala 131:10:@9517.4]
  assign _T_8814 = 4'hd <= offsetQ_4; // @[LoadQueue.scala 131:81:@9520.4]
  assign _T_8815 = _T_6344 & _T_8814; // @[LoadQueue.scala 131:72:@9521.4]
  assign _T_8817 = offsetQ_4 < 4'hd; // @[LoadQueue.scala 132:33:@9522.4]
  assign _T_8820 = _T_8817 & _T_6353; // @[LoadQueue.scala 132:41:@9524.4]
  assign _T_8822 = _T_8820 == 1'h0; // @[LoadQueue.scala 132:9:@9525.4]
  assign storesToCheck_4_13 = _T_2356 ? _T_8815 : _T_8822; // @[LoadQueue.scala 131:10:@9526.4]
  assign _T_8828 = 4'he <= offsetQ_4; // @[LoadQueue.scala 131:81:@9529.4]
  assign _T_8829 = _T_6361 & _T_8828; // @[LoadQueue.scala 131:72:@9530.4]
  assign _T_8831 = offsetQ_4 < 4'he; // @[LoadQueue.scala 132:33:@9531.4]
  assign _T_8834 = _T_8831 & _T_6370; // @[LoadQueue.scala 132:41:@9533.4]
  assign _T_8836 = _T_8834 == 1'h0; // @[LoadQueue.scala 132:9:@9534.4]
  assign storesToCheck_4_14 = _T_2356 ? _T_8829 : _T_8836; // @[LoadQueue.scala 131:10:@9535.4]
  assign _T_8842 = 4'hf <= offsetQ_4; // @[LoadQueue.scala 131:81:@9538.4]
  assign storesToCheck_4_15 = _T_2356 ? _T_8842 : 1'h1; // @[LoadQueue.scala 131:10:@9544.4]
  assign storesToCheck_5_0 = _T_2386 ? _T_6123 : 1'h1; // @[LoadQueue.scala 131:10:@9586.4]
  assign _T_8892 = 4'h1 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9589.4]
  assign _T_8893 = _T_6140 & _T_8892; // @[LoadQueue.scala 131:72:@9590.4]
  assign _T_8895 = offsetQ_5 < 4'h1; // @[LoadQueue.scala 132:33:@9591.4]
  assign _T_8898 = _T_8895 & _T_6149; // @[LoadQueue.scala 132:41:@9593.4]
  assign _T_8900 = _T_8898 == 1'h0; // @[LoadQueue.scala 132:9:@9594.4]
  assign storesToCheck_5_1 = _T_2386 ? _T_8893 : _T_8900; // @[LoadQueue.scala 131:10:@9595.4]
  assign _T_8906 = 4'h2 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9598.4]
  assign _T_8907 = _T_6157 & _T_8906; // @[LoadQueue.scala 131:72:@9599.4]
  assign _T_8909 = offsetQ_5 < 4'h2; // @[LoadQueue.scala 132:33:@9600.4]
  assign _T_8912 = _T_8909 & _T_6166; // @[LoadQueue.scala 132:41:@9602.4]
  assign _T_8914 = _T_8912 == 1'h0; // @[LoadQueue.scala 132:9:@9603.4]
  assign storesToCheck_5_2 = _T_2386 ? _T_8907 : _T_8914; // @[LoadQueue.scala 131:10:@9604.4]
  assign _T_8920 = 4'h3 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9607.4]
  assign _T_8921 = _T_6174 & _T_8920; // @[LoadQueue.scala 131:72:@9608.4]
  assign _T_8923 = offsetQ_5 < 4'h3; // @[LoadQueue.scala 132:33:@9609.4]
  assign _T_8926 = _T_8923 & _T_6183; // @[LoadQueue.scala 132:41:@9611.4]
  assign _T_8928 = _T_8926 == 1'h0; // @[LoadQueue.scala 132:9:@9612.4]
  assign storesToCheck_5_3 = _T_2386 ? _T_8921 : _T_8928; // @[LoadQueue.scala 131:10:@9613.4]
  assign _T_8934 = 4'h4 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9616.4]
  assign _T_8935 = _T_6191 & _T_8934; // @[LoadQueue.scala 131:72:@9617.4]
  assign _T_8937 = offsetQ_5 < 4'h4; // @[LoadQueue.scala 132:33:@9618.4]
  assign _T_8940 = _T_8937 & _T_6200; // @[LoadQueue.scala 132:41:@9620.4]
  assign _T_8942 = _T_8940 == 1'h0; // @[LoadQueue.scala 132:9:@9621.4]
  assign storesToCheck_5_4 = _T_2386 ? _T_8935 : _T_8942; // @[LoadQueue.scala 131:10:@9622.4]
  assign _T_8948 = 4'h5 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9625.4]
  assign _T_8949 = _T_6208 & _T_8948; // @[LoadQueue.scala 131:72:@9626.4]
  assign _T_8951 = offsetQ_5 < 4'h5; // @[LoadQueue.scala 132:33:@9627.4]
  assign _T_8954 = _T_8951 & _T_6217; // @[LoadQueue.scala 132:41:@9629.4]
  assign _T_8956 = _T_8954 == 1'h0; // @[LoadQueue.scala 132:9:@9630.4]
  assign storesToCheck_5_5 = _T_2386 ? _T_8949 : _T_8956; // @[LoadQueue.scala 131:10:@9631.4]
  assign _T_8962 = 4'h6 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9634.4]
  assign _T_8963 = _T_6225 & _T_8962; // @[LoadQueue.scala 131:72:@9635.4]
  assign _T_8965 = offsetQ_5 < 4'h6; // @[LoadQueue.scala 132:33:@9636.4]
  assign _T_8968 = _T_8965 & _T_6234; // @[LoadQueue.scala 132:41:@9638.4]
  assign _T_8970 = _T_8968 == 1'h0; // @[LoadQueue.scala 132:9:@9639.4]
  assign storesToCheck_5_6 = _T_2386 ? _T_8963 : _T_8970; // @[LoadQueue.scala 131:10:@9640.4]
  assign _T_8976 = 4'h7 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9643.4]
  assign _T_8977 = _T_6242 & _T_8976; // @[LoadQueue.scala 131:72:@9644.4]
  assign _T_8979 = offsetQ_5 < 4'h7; // @[LoadQueue.scala 132:33:@9645.4]
  assign _T_8982 = _T_8979 & _T_6251; // @[LoadQueue.scala 132:41:@9647.4]
  assign _T_8984 = _T_8982 == 1'h0; // @[LoadQueue.scala 132:9:@9648.4]
  assign storesToCheck_5_7 = _T_2386 ? _T_8977 : _T_8984; // @[LoadQueue.scala 131:10:@9649.4]
  assign _T_8990 = 4'h8 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9652.4]
  assign _T_8991 = _T_6259 & _T_8990; // @[LoadQueue.scala 131:72:@9653.4]
  assign _T_8993 = offsetQ_5 < 4'h8; // @[LoadQueue.scala 132:33:@9654.4]
  assign _T_8996 = _T_8993 & _T_6268; // @[LoadQueue.scala 132:41:@9656.4]
  assign _T_8998 = _T_8996 == 1'h0; // @[LoadQueue.scala 132:9:@9657.4]
  assign storesToCheck_5_8 = _T_2386 ? _T_8991 : _T_8998; // @[LoadQueue.scala 131:10:@9658.4]
  assign _T_9004 = 4'h9 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9661.4]
  assign _T_9005 = _T_6276 & _T_9004; // @[LoadQueue.scala 131:72:@9662.4]
  assign _T_9007 = offsetQ_5 < 4'h9; // @[LoadQueue.scala 132:33:@9663.4]
  assign _T_9010 = _T_9007 & _T_6285; // @[LoadQueue.scala 132:41:@9665.4]
  assign _T_9012 = _T_9010 == 1'h0; // @[LoadQueue.scala 132:9:@9666.4]
  assign storesToCheck_5_9 = _T_2386 ? _T_9005 : _T_9012; // @[LoadQueue.scala 131:10:@9667.4]
  assign _T_9018 = 4'ha <= offsetQ_5; // @[LoadQueue.scala 131:81:@9670.4]
  assign _T_9019 = _T_6293 & _T_9018; // @[LoadQueue.scala 131:72:@9671.4]
  assign _T_9021 = offsetQ_5 < 4'ha; // @[LoadQueue.scala 132:33:@9672.4]
  assign _T_9024 = _T_9021 & _T_6302; // @[LoadQueue.scala 132:41:@9674.4]
  assign _T_9026 = _T_9024 == 1'h0; // @[LoadQueue.scala 132:9:@9675.4]
  assign storesToCheck_5_10 = _T_2386 ? _T_9019 : _T_9026; // @[LoadQueue.scala 131:10:@9676.4]
  assign _T_9032 = 4'hb <= offsetQ_5; // @[LoadQueue.scala 131:81:@9679.4]
  assign _T_9033 = _T_6310 & _T_9032; // @[LoadQueue.scala 131:72:@9680.4]
  assign _T_9035 = offsetQ_5 < 4'hb; // @[LoadQueue.scala 132:33:@9681.4]
  assign _T_9038 = _T_9035 & _T_6319; // @[LoadQueue.scala 132:41:@9683.4]
  assign _T_9040 = _T_9038 == 1'h0; // @[LoadQueue.scala 132:9:@9684.4]
  assign storesToCheck_5_11 = _T_2386 ? _T_9033 : _T_9040; // @[LoadQueue.scala 131:10:@9685.4]
  assign _T_9046 = 4'hc <= offsetQ_5; // @[LoadQueue.scala 131:81:@9688.4]
  assign _T_9047 = _T_6327 & _T_9046; // @[LoadQueue.scala 131:72:@9689.4]
  assign _T_9049 = offsetQ_5 < 4'hc; // @[LoadQueue.scala 132:33:@9690.4]
  assign _T_9052 = _T_9049 & _T_6336; // @[LoadQueue.scala 132:41:@9692.4]
  assign _T_9054 = _T_9052 == 1'h0; // @[LoadQueue.scala 132:9:@9693.4]
  assign storesToCheck_5_12 = _T_2386 ? _T_9047 : _T_9054; // @[LoadQueue.scala 131:10:@9694.4]
  assign _T_9060 = 4'hd <= offsetQ_5; // @[LoadQueue.scala 131:81:@9697.4]
  assign _T_9061 = _T_6344 & _T_9060; // @[LoadQueue.scala 131:72:@9698.4]
  assign _T_9063 = offsetQ_5 < 4'hd; // @[LoadQueue.scala 132:33:@9699.4]
  assign _T_9066 = _T_9063 & _T_6353; // @[LoadQueue.scala 132:41:@9701.4]
  assign _T_9068 = _T_9066 == 1'h0; // @[LoadQueue.scala 132:9:@9702.4]
  assign storesToCheck_5_13 = _T_2386 ? _T_9061 : _T_9068; // @[LoadQueue.scala 131:10:@9703.4]
  assign _T_9074 = 4'he <= offsetQ_5; // @[LoadQueue.scala 131:81:@9706.4]
  assign _T_9075 = _T_6361 & _T_9074; // @[LoadQueue.scala 131:72:@9707.4]
  assign _T_9077 = offsetQ_5 < 4'he; // @[LoadQueue.scala 132:33:@9708.4]
  assign _T_9080 = _T_9077 & _T_6370; // @[LoadQueue.scala 132:41:@9710.4]
  assign _T_9082 = _T_9080 == 1'h0; // @[LoadQueue.scala 132:9:@9711.4]
  assign storesToCheck_5_14 = _T_2386 ? _T_9075 : _T_9082; // @[LoadQueue.scala 131:10:@9712.4]
  assign _T_9088 = 4'hf <= offsetQ_5; // @[LoadQueue.scala 131:81:@9715.4]
  assign storesToCheck_5_15 = _T_2386 ? _T_9088 : 1'h1; // @[LoadQueue.scala 131:10:@9721.4]
  assign storesToCheck_6_0 = _T_2416 ? _T_6123 : 1'h1; // @[LoadQueue.scala 131:10:@9763.4]
  assign _T_9138 = 4'h1 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9766.4]
  assign _T_9139 = _T_6140 & _T_9138; // @[LoadQueue.scala 131:72:@9767.4]
  assign _T_9141 = offsetQ_6 < 4'h1; // @[LoadQueue.scala 132:33:@9768.4]
  assign _T_9144 = _T_9141 & _T_6149; // @[LoadQueue.scala 132:41:@9770.4]
  assign _T_9146 = _T_9144 == 1'h0; // @[LoadQueue.scala 132:9:@9771.4]
  assign storesToCheck_6_1 = _T_2416 ? _T_9139 : _T_9146; // @[LoadQueue.scala 131:10:@9772.4]
  assign _T_9152 = 4'h2 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9775.4]
  assign _T_9153 = _T_6157 & _T_9152; // @[LoadQueue.scala 131:72:@9776.4]
  assign _T_9155 = offsetQ_6 < 4'h2; // @[LoadQueue.scala 132:33:@9777.4]
  assign _T_9158 = _T_9155 & _T_6166; // @[LoadQueue.scala 132:41:@9779.4]
  assign _T_9160 = _T_9158 == 1'h0; // @[LoadQueue.scala 132:9:@9780.4]
  assign storesToCheck_6_2 = _T_2416 ? _T_9153 : _T_9160; // @[LoadQueue.scala 131:10:@9781.4]
  assign _T_9166 = 4'h3 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9784.4]
  assign _T_9167 = _T_6174 & _T_9166; // @[LoadQueue.scala 131:72:@9785.4]
  assign _T_9169 = offsetQ_6 < 4'h3; // @[LoadQueue.scala 132:33:@9786.4]
  assign _T_9172 = _T_9169 & _T_6183; // @[LoadQueue.scala 132:41:@9788.4]
  assign _T_9174 = _T_9172 == 1'h0; // @[LoadQueue.scala 132:9:@9789.4]
  assign storesToCheck_6_3 = _T_2416 ? _T_9167 : _T_9174; // @[LoadQueue.scala 131:10:@9790.4]
  assign _T_9180 = 4'h4 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9793.4]
  assign _T_9181 = _T_6191 & _T_9180; // @[LoadQueue.scala 131:72:@9794.4]
  assign _T_9183 = offsetQ_6 < 4'h4; // @[LoadQueue.scala 132:33:@9795.4]
  assign _T_9186 = _T_9183 & _T_6200; // @[LoadQueue.scala 132:41:@9797.4]
  assign _T_9188 = _T_9186 == 1'h0; // @[LoadQueue.scala 132:9:@9798.4]
  assign storesToCheck_6_4 = _T_2416 ? _T_9181 : _T_9188; // @[LoadQueue.scala 131:10:@9799.4]
  assign _T_9194 = 4'h5 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9802.4]
  assign _T_9195 = _T_6208 & _T_9194; // @[LoadQueue.scala 131:72:@9803.4]
  assign _T_9197 = offsetQ_6 < 4'h5; // @[LoadQueue.scala 132:33:@9804.4]
  assign _T_9200 = _T_9197 & _T_6217; // @[LoadQueue.scala 132:41:@9806.4]
  assign _T_9202 = _T_9200 == 1'h0; // @[LoadQueue.scala 132:9:@9807.4]
  assign storesToCheck_6_5 = _T_2416 ? _T_9195 : _T_9202; // @[LoadQueue.scala 131:10:@9808.4]
  assign _T_9208 = 4'h6 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9811.4]
  assign _T_9209 = _T_6225 & _T_9208; // @[LoadQueue.scala 131:72:@9812.4]
  assign _T_9211 = offsetQ_6 < 4'h6; // @[LoadQueue.scala 132:33:@9813.4]
  assign _T_9214 = _T_9211 & _T_6234; // @[LoadQueue.scala 132:41:@9815.4]
  assign _T_9216 = _T_9214 == 1'h0; // @[LoadQueue.scala 132:9:@9816.4]
  assign storesToCheck_6_6 = _T_2416 ? _T_9209 : _T_9216; // @[LoadQueue.scala 131:10:@9817.4]
  assign _T_9222 = 4'h7 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9820.4]
  assign _T_9223 = _T_6242 & _T_9222; // @[LoadQueue.scala 131:72:@9821.4]
  assign _T_9225 = offsetQ_6 < 4'h7; // @[LoadQueue.scala 132:33:@9822.4]
  assign _T_9228 = _T_9225 & _T_6251; // @[LoadQueue.scala 132:41:@9824.4]
  assign _T_9230 = _T_9228 == 1'h0; // @[LoadQueue.scala 132:9:@9825.4]
  assign storesToCheck_6_7 = _T_2416 ? _T_9223 : _T_9230; // @[LoadQueue.scala 131:10:@9826.4]
  assign _T_9236 = 4'h8 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9829.4]
  assign _T_9237 = _T_6259 & _T_9236; // @[LoadQueue.scala 131:72:@9830.4]
  assign _T_9239 = offsetQ_6 < 4'h8; // @[LoadQueue.scala 132:33:@9831.4]
  assign _T_9242 = _T_9239 & _T_6268; // @[LoadQueue.scala 132:41:@9833.4]
  assign _T_9244 = _T_9242 == 1'h0; // @[LoadQueue.scala 132:9:@9834.4]
  assign storesToCheck_6_8 = _T_2416 ? _T_9237 : _T_9244; // @[LoadQueue.scala 131:10:@9835.4]
  assign _T_9250 = 4'h9 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9838.4]
  assign _T_9251 = _T_6276 & _T_9250; // @[LoadQueue.scala 131:72:@9839.4]
  assign _T_9253 = offsetQ_6 < 4'h9; // @[LoadQueue.scala 132:33:@9840.4]
  assign _T_9256 = _T_9253 & _T_6285; // @[LoadQueue.scala 132:41:@9842.4]
  assign _T_9258 = _T_9256 == 1'h0; // @[LoadQueue.scala 132:9:@9843.4]
  assign storesToCheck_6_9 = _T_2416 ? _T_9251 : _T_9258; // @[LoadQueue.scala 131:10:@9844.4]
  assign _T_9264 = 4'ha <= offsetQ_6; // @[LoadQueue.scala 131:81:@9847.4]
  assign _T_9265 = _T_6293 & _T_9264; // @[LoadQueue.scala 131:72:@9848.4]
  assign _T_9267 = offsetQ_6 < 4'ha; // @[LoadQueue.scala 132:33:@9849.4]
  assign _T_9270 = _T_9267 & _T_6302; // @[LoadQueue.scala 132:41:@9851.4]
  assign _T_9272 = _T_9270 == 1'h0; // @[LoadQueue.scala 132:9:@9852.4]
  assign storesToCheck_6_10 = _T_2416 ? _T_9265 : _T_9272; // @[LoadQueue.scala 131:10:@9853.4]
  assign _T_9278 = 4'hb <= offsetQ_6; // @[LoadQueue.scala 131:81:@9856.4]
  assign _T_9279 = _T_6310 & _T_9278; // @[LoadQueue.scala 131:72:@9857.4]
  assign _T_9281 = offsetQ_6 < 4'hb; // @[LoadQueue.scala 132:33:@9858.4]
  assign _T_9284 = _T_9281 & _T_6319; // @[LoadQueue.scala 132:41:@9860.4]
  assign _T_9286 = _T_9284 == 1'h0; // @[LoadQueue.scala 132:9:@9861.4]
  assign storesToCheck_6_11 = _T_2416 ? _T_9279 : _T_9286; // @[LoadQueue.scala 131:10:@9862.4]
  assign _T_9292 = 4'hc <= offsetQ_6; // @[LoadQueue.scala 131:81:@9865.4]
  assign _T_9293 = _T_6327 & _T_9292; // @[LoadQueue.scala 131:72:@9866.4]
  assign _T_9295 = offsetQ_6 < 4'hc; // @[LoadQueue.scala 132:33:@9867.4]
  assign _T_9298 = _T_9295 & _T_6336; // @[LoadQueue.scala 132:41:@9869.4]
  assign _T_9300 = _T_9298 == 1'h0; // @[LoadQueue.scala 132:9:@9870.4]
  assign storesToCheck_6_12 = _T_2416 ? _T_9293 : _T_9300; // @[LoadQueue.scala 131:10:@9871.4]
  assign _T_9306 = 4'hd <= offsetQ_6; // @[LoadQueue.scala 131:81:@9874.4]
  assign _T_9307 = _T_6344 & _T_9306; // @[LoadQueue.scala 131:72:@9875.4]
  assign _T_9309 = offsetQ_6 < 4'hd; // @[LoadQueue.scala 132:33:@9876.4]
  assign _T_9312 = _T_9309 & _T_6353; // @[LoadQueue.scala 132:41:@9878.4]
  assign _T_9314 = _T_9312 == 1'h0; // @[LoadQueue.scala 132:9:@9879.4]
  assign storesToCheck_6_13 = _T_2416 ? _T_9307 : _T_9314; // @[LoadQueue.scala 131:10:@9880.4]
  assign _T_9320 = 4'he <= offsetQ_6; // @[LoadQueue.scala 131:81:@9883.4]
  assign _T_9321 = _T_6361 & _T_9320; // @[LoadQueue.scala 131:72:@9884.4]
  assign _T_9323 = offsetQ_6 < 4'he; // @[LoadQueue.scala 132:33:@9885.4]
  assign _T_9326 = _T_9323 & _T_6370; // @[LoadQueue.scala 132:41:@9887.4]
  assign _T_9328 = _T_9326 == 1'h0; // @[LoadQueue.scala 132:9:@9888.4]
  assign storesToCheck_6_14 = _T_2416 ? _T_9321 : _T_9328; // @[LoadQueue.scala 131:10:@9889.4]
  assign _T_9334 = 4'hf <= offsetQ_6; // @[LoadQueue.scala 131:81:@9892.4]
  assign storesToCheck_6_15 = _T_2416 ? _T_9334 : 1'h1; // @[LoadQueue.scala 131:10:@9898.4]
  assign storesToCheck_7_0 = _T_2446 ? _T_6123 : 1'h1; // @[LoadQueue.scala 131:10:@9940.4]
  assign _T_9384 = 4'h1 <= offsetQ_7; // @[LoadQueue.scala 131:81:@9943.4]
  assign _T_9385 = _T_6140 & _T_9384; // @[LoadQueue.scala 131:72:@9944.4]
  assign _T_9387 = offsetQ_7 < 4'h1; // @[LoadQueue.scala 132:33:@9945.4]
  assign _T_9390 = _T_9387 & _T_6149; // @[LoadQueue.scala 132:41:@9947.4]
  assign _T_9392 = _T_9390 == 1'h0; // @[LoadQueue.scala 132:9:@9948.4]
  assign storesToCheck_7_1 = _T_2446 ? _T_9385 : _T_9392; // @[LoadQueue.scala 131:10:@9949.4]
  assign _T_9398 = 4'h2 <= offsetQ_7; // @[LoadQueue.scala 131:81:@9952.4]
  assign _T_9399 = _T_6157 & _T_9398; // @[LoadQueue.scala 131:72:@9953.4]
  assign _T_9401 = offsetQ_7 < 4'h2; // @[LoadQueue.scala 132:33:@9954.4]
  assign _T_9404 = _T_9401 & _T_6166; // @[LoadQueue.scala 132:41:@9956.4]
  assign _T_9406 = _T_9404 == 1'h0; // @[LoadQueue.scala 132:9:@9957.4]
  assign storesToCheck_7_2 = _T_2446 ? _T_9399 : _T_9406; // @[LoadQueue.scala 131:10:@9958.4]
  assign _T_9412 = 4'h3 <= offsetQ_7; // @[LoadQueue.scala 131:81:@9961.4]
  assign _T_9413 = _T_6174 & _T_9412; // @[LoadQueue.scala 131:72:@9962.4]
  assign _T_9415 = offsetQ_7 < 4'h3; // @[LoadQueue.scala 132:33:@9963.4]
  assign _T_9418 = _T_9415 & _T_6183; // @[LoadQueue.scala 132:41:@9965.4]
  assign _T_9420 = _T_9418 == 1'h0; // @[LoadQueue.scala 132:9:@9966.4]
  assign storesToCheck_7_3 = _T_2446 ? _T_9413 : _T_9420; // @[LoadQueue.scala 131:10:@9967.4]
  assign _T_9426 = 4'h4 <= offsetQ_7; // @[LoadQueue.scala 131:81:@9970.4]
  assign _T_9427 = _T_6191 & _T_9426; // @[LoadQueue.scala 131:72:@9971.4]
  assign _T_9429 = offsetQ_7 < 4'h4; // @[LoadQueue.scala 132:33:@9972.4]
  assign _T_9432 = _T_9429 & _T_6200; // @[LoadQueue.scala 132:41:@9974.4]
  assign _T_9434 = _T_9432 == 1'h0; // @[LoadQueue.scala 132:9:@9975.4]
  assign storesToCheck_7_4 = _T_2446 ? _T_9427 : _T_9434; // @[LoadQueue.scala 131:10:@9976.4]
  assign _T_9440 = 4'h5 <= offsetQ_7; // @[LoadQueue.scala 131:81:@9979.4]
  assign _T_9441 = _T_6208 & _T_9440; // @[LoadQueue.scala 131:72:@9980.4]
  assign _T_9443 = offsetQ_7 < 4'h5; // @[LoadQueue.scala 132:33:@9981.4]
  assign _T_9446 = _T_9443 & _T_6217; // @[LoadQueue.scala 132:41:@9983.4]
  assign _T_9448 = _T_9446 == 1'h0; // @[LoadQueue.scala 132:9:@9984.4]
  assign storesToCheck_7_5 = _T_2446 ? _T_9441 : _T_9448; // @[LoadQueue.scala 131:10:@9985.4]
  assign _T_9454 = 4'h6 <= offsetQ_7; // @[LoadQueue.scala 131:81:@9988.4]
  assign _T_9455 = _T_6225 & _T_9454; // @[LoadQueue.scala 131:72:@9989.4]
  assign _T_9457 = offsetQ_7 < 4'h6; // @[LoadQueue.scala 132:33:@9990.4]
  assign _T_9460 = _T_9457 & _T_6234; // @[LoadQueue.scala 132:41:@9992.4]
  assign _T_9462 = _T_9460 == 1'h0; // @[LoadQueue.scala 132:9:@9993.4]
  assign storesToCheck_7_6 = _T_2446 ? _T_9455 : _T_9462; // @[LoadQueue.scala 131:10:@9994.4]
  assign _T_9468 = 4'h7 <= offsetQ_7; // @[LoadQueue.scala 131:81:@9997.4]
  assign _T_9469 = _T_6242 & _T_9468; // @[LoadQueue.scala 131:72:@9998.4]
  assign _T_9471 = offsetQ_7 < 4'h7; // @[LoadQueue.scala 132:33:@9999.4]
  assign _T_9474 = _T_9471 & _T_6251; // @[LoadQueue.scala 132:41:@10001.4]
  assign _T_9476 = _T_9474 == 1'h0; // @[LoadQueue.scala 132:9:@10002.4]
  assign storesToCheck_7_7 = _T_2446 ? _T_9469 : _T_9476; // @[LoadQueue.scala 131:10:@10003.4]
  assign _T_9482 = 4'h8 <= offsetQ_7; // @[LoadQueue.scala 131:81:@10006.4]
  assign _T_9483 = _T_6259 & _T_9482; // @[LoadQueue.scala 131:72:@10007.4]
  assign _T_9485 = offsetQ_7 < 4'h8; // @[LoadQueue.scala 132:33:@10008.4]
  assign _T_9488 = _T_9485 & _T_6268; // @[LoadQueue.scala 132:41:@10010.4]
  assign _T_9490 = _T_9488 == 1'h0; // @[LoadQueue.scala 132:9:@10011.4]
  assign storesToCheck_7_8 = _T_2446 ? _T_9483 : _T_9490; // @[LoadQueue.scala 131:10:@10012.4]
  assign _T_9496 = 4'h9 <= offsetQ_7; // @[LoadQueue.scala 131:81:@10015.4]
  assign _T_9497 = _T_6276 & _T_9496; // @[LoadQueue.scala 131:72:@10016.4]
  assign _T_9499 = offsetQ_7 < 4'h9; // @[LoadQueue.scala 132:33:@10017.4]
  assign _T_9502 = _T_9499 & _T_6285; // @[LoadQueue.scala 132:41:@10019.4]
  assign _T_9504 = _T_9502 == 1'h0; // @[LoadQueue.scala 132:9:@10020.4]
  assign storesToCheck_7_9 = _T_2446 ? _T_9497 : _T_9504; // @[LoadQueue.scala 131:10:@10021.4]
  assign _T_9510 = 4'ha <= offsetQ_7; // @[LoadQueue.scala 131:81:@10024.4]
  assign _T_9511 = _T_6293 & _T_9510; // @[LoadQueue.scala 131:72:@10025.4]
  assign _T_9513 = offsetQ_7 < 4'ha; // @[LoadQueue.scala 132:33:@10026.4]
  assign _T_9516 = _T_9513 & _T_6302; // @[LoadQueue.scala 132:41:@10028.4]
  assign _T_9518 = _T_9516 == 1'h0; // @[LoadQueue.scala 132:9:@10029.4]
  assign storesToCheck_7_10 = _T_2446 ? _T_9511 : _T_9518; // @[LoadQueue.scala 131:10:@10030.4]
  assign _T_9524 = 4'hb <= offsetQ_7; // @[LoadQueue.scala 131:81:@10033.4]
  assign _T_9525 = _T_6310 & _T_9524; // @[LoadQueue.scala 131:72:@10034.4]
  assign _T_9527 = offsetQ_7 < 4'hb; // @[LoadQueue.scala 132:33:@10035.4]
  assign _T_9530 = _T_9527 & _T_6319; // @[LoadQueue.scala 132:41:@10037.4]
  assign _T_9532 = _T_9530 == 1'h0; // @[LoadQueue.scala 132:9:@10038.4]
  assign storesToCheck_7_11 = _T_2446 ? _T_9525 : _T_9532; // @[LoadQueue.scala 131:10:@10039.4]
  assign _T_9538 = 4'hc <= offsetQ_7; // @[LoadQueue.scala 131:81:@10042.4]
  assign _T_9539 = _T_6327 & _T_9538; // @[LoadQueue.scala 131:72:@10043.4]
  assign _T_9541 = offsetQ_7 < 4'hc; // @[LoadQueue.scala 132:33:@10044.4]
  assign _T_9544 = _T_9541 & _T_6336; // @[LoadQueue.scala 132:41:@10046.4]
  assign _T_9546 = _T_9544 == 1'h0; // @[LoadQueue.scala 132:9:@10047.4]
  assign storesToCheck_7_12 = _T_2446 ? _T_9539 : _T_9546; // @[LoadQueue.scala 131:10:@10048.4]
  assign _T_9552 = 4'hd <= offsetQ_7; // @[LoadQueue.scala 131:81:@10051.4]
  assign _T_9553 = _T_6344 & _T_9552; // @[LoadQueue.scala 131:72:@10052.4]
  assign _T_9555 = offsetQ_7 < 4'hd; // @[LoadQueue.scala 132:33:@10053.4]
  assign _T_9558 = _T_9555 & _T_6353; // @[LoadQueue.scala 132:41:@10055.4]
  assign _T_9560 = _T_9558 == 1'h0; // @[LoadQueue.scala 132:9:@10056.4]
  assign storesToCheck_7_13 = _T_2446 ? _T_9553 : _T_9560; // @[LoadQueue.scala 131:10:@10057.4]
  assign _T_9566 = 4'he <= offsetQ_7; // @[LoadQueue.scala 131:81:@10060.4]
  assign _T_9567 = _T_6361 & _T_9566; // @[LoadQueue.scala 131:72:@10061.4]
  assign _T_9569 = offsetQ_7 < 4'he; // @[LoadQueue.scala 132:33:@10062.4]
  assign _T_9572 = _T_9569 & _T_6370; // @[LoadQueue.scala 132:41:@10064.4]
  assign _T_9574 = _T_9572 == 1'h0; // @[LoadQueue.scala 132:9:@10065.4]
  assign storesToCheck_7_14 = _T_2446 ? _T_9567 : _T_9574; // @[LoadQueue.scala 131:10:@10066.4]
  assign _T_9580 = 4'hf <= offsetQ_7; // @[LoadQueue.scala 131:81:@10069.4]
  assign storesToCheck_7_15 = _T_2446 ? _T_9580 : 1'h1; // @[LoadQueue.scala 131:10:@10075.4]
  assign storesToCheck_8_0 = _T_2476 ? _T_6123 : 1'h1; // @[LoadQueue.scala 131:10:@10117.4]
  assign _T_9630 = 4'h1 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10120.4]
  assign _T_9631 = _T_6140 & _T_9630; // @[LoadQueue.scala 131:72:@10121.4]
  assign _T_9633 = offsetQ_8 < 4'h1; // @[LoadQueue.scala 132:33:@10122.4]
  assign _T_9636 = _T_9633 & _T_6149; // @[LoadQueue.scala 132:41:@10124.4]
  assign _T_9638 = _T_9636 == 1'h0; // @[LoadQueue.scala 132:9:@10125.4]
  assign storesToCheck_8_1 = _T_2476 ? _T_9631 : _T_9638; // @[LoadQueue.scala 131:10:@10126.4]
  assign _T_9644 = 4'h2 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10129.4]
  assign _T_9645 = _T_6157 & _T_9644; // @[LoadQueue.scala 131:72:@10130.4]
  assign _T_9647 = offsetQ_8 < 4'h2; // @[LoadQueue.scala 132:33:@10131.4]
  assign _T_9650 = _T_9647 & _T_6166; // @[LoadQueue.scala 132:41:@10133.4]
  assign _T_9652 = _T_9650 == 1'h0; // @[LoadQueue.scala 132:9:@10134.4]
  assign storesToCheck_8_2 = _T_2476 ? _T_9645 : _T_9652; // @[LoadQueue.scala 131:10:@10135.4]
  assign _T_9658 = 4'h3 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10138.4]
  assign _T_9659 = _T_6174 & _T_9658; // @[LoadQueue.scala 131:72:@10139.4]
  assign _T_9661 = offsetQ_8 < 4'h3; // @[LoadQueue.scala 132:33:@10140.4]
  assign _T_9664 = _T_9661 & _T_6183; // @[LoadQueue.scala 132:41:@10142.4]
  assign _T_9666 = _T_9664 == 1'h0; // @[LoadQueue.scala 132:9:@10143.4]
  assign storesToCheck_8_3 = _T_2476 ? _T_9659 : _T_9666; // @[LoadQueue.scala 131:10:@10144.4]
  assign _T_9672 = 4'h4 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10147.4]
  assign _T_9673 = _T_6191 & _T_9672; // @[LoadQueue.scala 131:72:@10148.4]
  assign _T_9675 = offsetQ_8 < 4'h4; // @[LoadQueue.scala 132:33:@10149.4]
  assign _T_9678 = _T_9675 & _T_6200; // @[LoadQueue.scala 132:41:@10151.4]
  assign _T_9680 = _T_9678 == 1'h0; // @[LoadQueue.scala 132:9:@10152.4]
  assign storesToCheck_8_4 = _T_2476 ? _T_9673 : _T_9680; // @[LoadQueue.scala 131:10:@10153.4]
  assign _T_9686 = 4'h5 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10156.4]
  assign _T_9687 = _T_6208 & _T_9686; // @[LoadQueue.scala 131:72:@10157.4]
  assign _T_9689 = offsetQ_8 < 4'h5; // @[LoadQueue.scala 132:33:@10158.4]
  assign _T_9692 = _T_9689 & _T_6217; // @[LoadQueue.scala 132:41:@10160.4]
  assign _T_9694 = _T_9692 == 1'h0; // @[LoadQueue.scala 132:9:@10161.4]
  assign storesToCheck_8_5 = _T_2476 ? _T_9687 : _T_9694; // @[LoadQueue.scala 131:10:@10162.4]
  assign _T_9700 = 4'h6 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10165.4]
  assign _T_9701 = _T_6225 & _T_9700; // @[LoadQueue.scala 131:72:@10166.4]
  assign _T_9703 = offsetQ_8 < 4'h6; // @[LoadQueue.scala 132:33:@10167.4]
  assign _T_9706 = _T_9703 & _T_6234; // @[LoadQueue.scala 132:41:@10169.4]
  assign _T_9708 = _T_9706 == 1'h0; // @[LoadQueue.scala 132:9:@10170.4]
  assign storesToCheck_8_6 = _T_2476 ? _T_9701 : _T_9708; // @[LoadQueue.scala 131:10:@10171.4]
  assign _T_9714 = 4'h7 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10174.4]
  assign _T_9715 = _T_6242 & _T_9714; // @[LoadQueue.scala 131:72:@10175.4]
  assign _T_9717 = offsetQ_8 < 4'h7; // @[LoadQueue.scala 132:33:@10176.4]
  assign _T_9720 = _T_9717 & _T_6251; // @[LoadQueue.scala 132:41:@10178.4]
  assign _T_9722 = _T_9720 == 1'h0; // @[LoadQueue.scala 132:9:@10179.4]
  assign storesToCheck_8_7 = _T_2476 ? _T_9715 : _T_9722; // @[LoadQueue.scala 131:10:@10180.4]
  assign _T_9728 = 4'h8 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10183.4]
  assign _T_9729 = _T_6259 & _T_9728; // @[LoadQueue.scala 131:72:@10184.4]
  assign _T_9731 = offsetQ_8 < 4'h8; // @[LoadQueue.scala 132:33:@10185.4]
  assign _T_9734 = _T_9731 & _T_6268; // @[LoadQueue.scala 132:41:@10187.4]
  assign _T_9736 = _T_9734 == 1'h0; // @[LoadQueue.scala 132:9:@10188.4]
  assign storesToCheck_8_8 = _T_2476 ? _T_9729 : _T_9736; // @[LoadQueue.scala 131:10:@10189.4]
  assign _T_9742 = 4'h9 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10192.4]
  assign _T_9743 = _T_6276 & _T_9742; // @[LoadQueue.scala 131:72:@10193.4]
  assign _T_9745 = offsetQ_8 < 4'h9; // @[LoadQueue.scala 132:33:@10194.4]
  assign _T_9748 = _T_9745 & _T_6285; // @[LoadQueue.scala 132:41:@10196.4]
  assign _T_9750 = _T_9748 == 1'h0; // @[LoadQueue.scala 132:9:@10197.4]
  assign storesToCheck_8_9 = _T_2476 ? _T_9743 : _T_9750; // @[LoadQueue.scala 131:10:@10198.4]
  assign _T_9756 = 4'ha <= offsetQ_8; // @[LoadQueue.scala 131:81:@10201.4]
  assign _T_9757 = _T_6293 & _T_9756; // @[LoadQueue.scala 131:72:@10202.4]
  assign _T_9759 = offsetQ_8 < 4'ha; // @[LoadQueue.scala 132:33:@10203.4]
  assign _T_9762 = _T_9759 & _T_6302; // @[LoadQueue.scala 132:41:@10205.4]
  assign _T_9764 = _T_9762 == 1'h0; // @[LoadQueue.scala 132:9:@10206.4]
  assign storesToCheck_8_10 = _T_2476 ? _T_9757 : _T_9764; // @[LoadQueue.scala 131:10:@10207.4]
  assign _T_9770 = 4'hb <= offsetQ_8; // @[LoadQueue.scala 131:81:@10210.4]
  assign _T_9771 = _T_6310 & _T_9770; // @[LoadQueue.scala 131:72:@10211.4]
  assign _T_9773 = offsetQ_8 < 4'hb; // @[LoadQueue.scala 132:33:@10212.4]
  assign _T_9776 = _T_9773 & _T_6319; // @[LoadQueue.scala 132:41:@10214.4]
  assign _T_9778 = _T_9776 == 1'h0; // @[LoadQueue.scala 132:9:@10215.4]
  assign storesToCheck_8_11 = _T_2476 ? _T_9771 : _T_9778; // @[LoadQueue.scala 131:10:@10216.4]
  assign _T_9784 = 4'hc <= offsetQ_8; // @[LoadQueue.scala 131:81:@10219.4]
  assign _T_9785 = _T_6327 & _T_9784; // @[LoadQueue.scala 131:72:@10220.4]
  assign _T_9787 = offsetQ_8 < 4'hc; // @[LoadQueue.scala 132:33:@10221.4]
  assign _T_9790 = _T_9787 & _T_6336; // @[LoadQueue.scala 132:41:@10223.4]
  assign _T_9792 = _T_9790 == 1'h0; // @[LoadQueue.scala 132:9:@10224.4]
  assign storesToCheck_8_12 = _T_2476 ? _T_9785 : _T_9792; // @[LoadQueue.scala 131:10:@10225.4]
  assign _T_9798 = 4'hd <= offsetQ_8; // @[LoadQueue.scala 131:81:@10228.4]
  assign _T_9799 = _T_6344 & _T_9798; // @[LoadQueue.scala 131:72:@10229.4]
  assign _T_9801 = offsetQ_8 < 4'hd; // @[LoadQueue.scala 132:33:@10230.4]
  assign _T_9804 = _T_9801 & _T_6353; // @[LoadQueue.scala 132:41:@10232.4]
  assign _T_9806 = _T_9804 == 1'h0; // @[LoadQueue.scala 132:9:@10233.4]
  assign storesToCheck_8_13 = _T_2476 ? _T_9799 : _T_9806; // @[LoadQueue.scala 131:10:@10234.4]
  assign _T_9812 = 4'he <= offsetQ_8; // @[LoadQueue.scala 131:81:@10237.4]
  assign _T_9813 = _T_6361 & _T_9812; // @[LoadQueue.scala 131:72:@10238.4]
  assign _T_9815 = offsetQ_8 < 4'he; // @[LoadQueue.scala 132:33:@10239.4]
  assign _T_9818 = _T_9815 & _T_6370; // @[LoadQueue.scala 132:41:@10241.4]
  assign _T_9820 = _T_9818 == 1'h0; // @[LoadQueue.scala 132:9:@10242.4]
  assign storesToCheck_8_14 = _T_2476 ? _T_9813 : _T_9820; // @[LoadQueue.scala 131:10:@10243.4]
  assign _T_9826 = 4'hf <= offsetQ_8; // @[LoadQueue.scala 131:81:@10246.4]
  assign storesToCheck_8_15 = _T_2476 ? _T_9826 : 1'h1; // @[LoadQueue.scala 131:10:@10252.4]
  assign storesToCheck_9_0 = _T_2506 ? _T_6123 : 1'h1; // @[LoadQueue.scala 131:10:@10294.4]
  assign _T_9876 = 4'h1 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10297.4]
  assign _T_9877 = _T_6140 & _T_9876; // @[LoadQueue.scala 131:72:@10298.4]
  assign _T_9879 = offsetQ_9 < 4'h1; // @[LoadQueue.scala 132:33:@10299.4]
  assign _T_9882 = _T_9879 & _T_6149; // @[LoadQueue.scala 132:41:@10301.4]
  assign _T_9884 = _T_9882 == 1'h0; // @[LoadQueue.scala 132:9:@10302.4]
  assign storesToCheck_9_1 = _T_2506 ? _T_9877 : _T_9884; // @[LoadQueue.scala 131:10:@10303.4]
  assign _T_9890 = 4'h2 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10306.4]
  assign _T_9891 = _T_6157 & _T_9890; // @[LoadQueue.scala 131:72:@10307.4]
  assign _T_9893 = offsetQ_9 < 4'h2; // @[LoadQueue.scala 132:33:@10308.4]
  assign _T_9896 = _T_9893 & _T_6166; // @[LoadQueue.scala 132:41:@10310.4]
  assign _T_9898 = _T_9896 == 1'h0; // @[LoadQueue.scala 132:9:@10311.4]
  assign storesToCheck_9_2 = _T_2506 ? _T_9891 : _T_9898; // @[LoadQueue.scala 131:10:@10312.4]
  assign _T_9904 = 4'h3 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10315.4]
  assign _T_9905 = _T_6174 & _T_9904; // @[LoadQueue.scala 131:72:@10316.4]
  assign _T_9907 = offsetQ_9 < 4'h3; // @[LoadQueue.scala 132:33:@10317.4]
  assign _T_9910 = _T_9907 & _T_6183; // @[LoadQueue.scala 132:41:@10319.4]
  assign _T_9912 = _T_9910 == 1'h0; // @[LoadQueue.scala 132:9:@10320.4]
  assign storesToCheck_9_3 = _T_2506 ? _T_9905 : _T_9912; // @[LoadQueue.scala 131:10:@10321.4]
  assign _T_9918 = 4'h4 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10324.4]
  assign _T_9919 = _T_6191 & _T_9918; // @[LoadQueue.scala 131:72:@10325.4]
  assign _T_9921 = offsetQ_9 < 4'h4; // @[LoadQueue.scala 132:33:@10326.4]
  assign _T_9924 = _T_9921 & _T_6200; // @[LoadQueue.scala 132:41:@10328.4]
  assign _T_9926 = _T_9924 == 1'h0; // @[LoadQueue.scala 132:9:@10329.4]
  assign storesToCheck_9_4 = _T_2506 ? _T_9919 : _T_9926; // @[LoadQueue.scala 131:10:@10330.4]
  assign _T_9932 = 4'h5 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10333.4]
  assign _T_9933 = _T_6208 & _T_9932; // @[LoadQueue.scala 131:72:@10334.4]
  assign _T_9935 = offsetQ_9 < 4'h5; // @[LoadQueue.scala 132:33:@10335.4]
  assign _T_9938 = _T_9935 & _T_6217; // @[LoadQueue.scala 132:41:@10337.4]
  assign _T_9940 = _T_9938 == 1'h0; // @[LoadQueue.scala 132:9:@10338.4]
  assign storesToCheck_9_5 = _T_2506 ? _T_9933 : _T_9940; // @[LoadQueue.scala 131:10:@10339.4]
  assign _T_9946 = 4'h6 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10342.4]
  assign _T_9947 = _T_6225 & _T_9946; // @[LoadQueue.scala 131:72:@10343.4]
  assign _T_9949 = offsetQ_9 < 4'h6; // @[LoadQueue.scala 132:33:@10344.4]
  assign _T_9952 = _T_9949 & _T_6234; // @[LoadQueue.scala 132:41:@10346.4]
  assign _T_9954 = _T_9952 == 1'h0; // @[LoadQueue.scala 132:9:@10347.4]
  assign storesToCheck_9_6 = _T_2506 ? _T_9947 : _T_9954; // @[LoadQueue.scala 131:10:@10348.4]
  assign _T_9960 = 4'h7 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10351.4]
  assign _T_9961 = _T_6242 & _T_9960; // @[LoadQueue.scala 131:72:@10352.4]
  assign _T_9963 = offsetQ_9 < 4'h7; // @[LoadQueue.scala 132:33:@10353.4]
  assign _T_9966 = _T_9963 & _T_6251; // @[LoadQueue.scala 132:41:@10355.4]
  assign _T_9968 = _T_9966 == 1'h0; // @[LoadQueue.scala 132:9:@10356.4]
  assign storesToCheck_9_7 = _T_2506 ? _T_9961 : _T_9968; // @[LoadQueue.scala 131:10:@10357.4]
  assign _T_9974 = 4'h8 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10360.4]
  assign _T_9975 = _T_6259 & _T_9974; // @[LoadQueue.scala 131:72:@10361.4]
  assign _T_9977 = offsetQ_9 < 4'h8; // @[LoadQueue.scala 132:33:@10362.4]
  assign _T_9980 = _T_9977 & _T_6268; // @[LoadQueue.scala 132:41:@10364.4]
  assign _T_9982 = _T_9980 == 1'h0; // @[LoadQueue.scala 132:9:@10365.4]
  assign storesToCheck_9_8 = _T_2506 ? _T_9975 : _T_9982; // @[LoadQueue.scala 131:10:@10366.4]
  assign _T_9988 = 4'h9 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10369.4]
  assign _T_9989 = _T_6276 & _T_9988; // @[LoadQueue.scala 131:72:@10370.4]
  assign _T_9991 = offsetQ_9 < 4'h9; // @[LoadQueue.scala 132:33:@10371.4]
  assign _T_9994 = _T_9991 & _T_6285; // @[LoadQueue.scala 132:41:@10373.4]
  assign _T_9996 = _T_9994 == 1'h0; // @[LoadQueue.scala 132:9:@10374.4]
  assign storesToCheck_9_9 = _T_2506 ? _T_9989 : _T_9996; // @[LoadQueue.scala 131:10:@10375.4]
  assign _T_10002 = 4'ha <= offsetQ_9; // @[LoadQueue.scala 131:81:@10378.4]
  assign _T_10003 = _T_6293 & _T_10002; // @[LoadQueue.scala 131:72:@10379.4]
  assign _T_10005 = offsetQ_9 < 4'ha; // @[LoadQueue.scala 132:33:@10380.4]
  assign _T_10008 = _T_10005 & _T_6302; // @[LoadQueue.scala 132:41:@10382.4]
  assign _T_10010 = _T_10008 == 1'h0; // @[LoadQueue.scala 132:9:@10383.4]
  assign storesToCheck_9_10 = _T_2506 ? _T_10003 : _T_10010; // @[LoadQueue.scala 131:10:@10384.4]
  assign _T_10016 = 4'hb <= offsetQ_9; // @[LoadQueue.scala 131:81:@10387.4]
  assign _T_10017 = _T_6310 & _T_10016; // @[LoadQueue.scala 131:72:@10388.4]
  assign _T_10019 = offsetQ_9 < 4'hb; // @[LoadQueue.scala 132:33:@10389.4]
  assign _T_10022 = _T_10019 & _T_6319; // @[LoadQueue.scala 132:41:@10391.4]
  assign _T_10024 = _T_10022 == 1'h0; // @[LoadQueue.scala 132:9:@10392.4]
  assign storesToCheck_9_11 = _T_2506 ? _T_10017 : _T_10024; // @[LoadQueue.scala 131:10:@10393.4]
  assign _T_10030 = 4'hc <= offsetQ_9; // @[LoadQueue.scala 131:81:@10396.4]
  assign _T_10031 = _T_6327 & _T_10030; // @[LoadQueue.scala 131:72:@10397.4]
  assign _T_10033 = offsetQ_9 < 4'hc; // @[LoadQueue.scala 132:33:@10398.4]
  assign _T_10036 = _T_10033 & _T_6336; // @[LoadQueue.scala 132:41:@10400.4]
  assign _T_10038 = _T_10036 == 1'h0; // @[LoadQueue.scala 132:9:@10401.4]
  assign storesToCheck_9_12 = _T_2506 ? _T_10031 : _T_10038; // @[LoadQueue.scala 131:10:@10402.4]
  assign _T_10044 = 4'hd <= offsetQ_9; // @[LoadQueue.scala 131:81:@10405.4]
  assign _T_10045 = _T_6344 & _T_10044; // @[LoadQueue.scala 131:72:@10406.4]
  assign _T_10047 = offsetQ_9 < 4'hd; // @[LoadQueue.scala 132:33:@10407.4]
  assign _T_10050 = _T_10047 & _T_6353; // @[LoadQueue.scala 132:41:@10409.4]
  assign _T_10052 = _T_10050 == 1'h0; // @[LoadQueue.scala 132:9:@10410.4]
  assign storesToCheck_9_13 = _T_2506 ? _T_10045 : _T_10052; // @[LoadQueue.scala 131:10:@10411.4]
  assign _T_10058 = 4'he <= offsetQ_9; // @[LoadQueue.scala 131:81:@10414.4]
  assign _T_10059 = _T_6361 & _T_10058; // @[LoadQueue.scala 131:72:@10415.4]
  assign _T_10061 = offsetQ_9 < 4'he; // @[LoadQueue.scala 132:33:@10416.4]
  assign _T_10064 = _T_10061 & _T_6370; // @[LoadQueue.scala 132:41:@10418.4]
  assign _T_10066 = _T_10064 == 1'h0; // @[LoadQueue.scala 132:9:@10419.4]
  assign storesToCheck_9_14 = _T_2506 ? _T_10059 : _T_10066; // @[LoadQueue.scala 131:10:@10420.4]
  assign _T_10072 = 4'hf <= offsetQ_9; // @[LoadQueue.scala 131:81:@10423.4]
  assign storesToCheck_9_15 = _T_2506 ? _T_10072 : 1'h1; // @[LoadQueue.scala 131:10:@10429.4]
  assign storesToCheck_10_0 = _T_2536 ? _T_6123 : 1'h1; // @[LoadQueue.scala 131:10:@10471.4]
  assign _T_10122 = 4'h1 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10474.4]
  assign _T_10123 = _T_6140 & _T_10122; // @[LoadQueue.scala 131:72:@10475.4]
  assign _T_10125 = offsetQ_10 < 4'h1; // @[LoadQueue.scala 132:33:@10476.4]
  assign _T_10128 = _T_10125 & _T_6149; // @[LoadQueue.scala 132:41:@10478.4]
  assign _T_10130 = _T_10128 == 1'h0; // @[LoadQueue.scala 132:9:@10479.4]
  assign storesToCheck_10_1 = _T_2536 ? _T_10123 : _T_10130; // @[LoadQueue.scala 131:10:@10480.4]
  assign _T_10136 = 4'h2 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10483.4]
  assign _T_10137 = _T_6157 & _T_10136; // @[LoadQueue.scala 131:72:@10484.4]
  assign _T_10139 = offsetQ_10 < 4'h2; // @[LoadQueue.scala 132:33:@10485.4]
  assign _T_10142 = _T_10139 & _T_6166; // @[LoadQueue.scala 132:41:@10487.4]
  assign _T_10144 = _T_10142 == 1'h0; // @[LoadQueue.scala 132:9:@10488.4]
  assign storesToCheck_10_2 = _T_2536 ? _T_10137 : _T_10144; // @[LoadQueue.scala 131:10:@10489.4]
  assign _T_10150 = 4'h3 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10492.4]
  assign _T_10151 = _T_6174 & _T_10150; // @[LoadQueue.scala 131:72:@10493.4]
  assign _T_10153 = offsetQ_10 < 4'h3; // @[LoadQueue.scala 132:33:@10494.4]
  assign _T_10156 = _T_10153 & _T_6183; // @[LoadQueue.scala 132:41:@10496.4]
  assign _T_10158 = _T_10156 == 1'h0; // @[LoadQueue.scala 132:9:@10497.4]
  assign storesToCheck_10_3 = _T_2536 ? _T_10151 : _T_10158; // @[LoadQueue.scala 131:10:@10498.4]
  assign _T_10164 = 4'h4 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10501.4]
  assign _T_10165 = _T_6191 & _T_10164; // @[LoadQueue.scala 131:72:@10502.4]
  assign _T_10167 = offsetQ_10 < 4'h4; // @[LoadQueue.scala 132:33:@10503.4]
  assign _T_10170 = _T_10167 & _T_6200; // @[LoadQueue.scala 132:41:@10505.4]
  assign _T_10172 = _T_10170 == 1'h0; // @[LoadQueue.scala 132:9:@10506.4]
  assign storesToCheck_10_4 = _T_2536 ? _T_10165 : _T_10172; // @[LoadQueue.scala 131:10:@10507.4]
  assign _T_10178 = 4'h5 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10510.4]
  assign _T_10179 = _T_6208 & _T_10178; // @[LoadQueue.scala 131:72:@10511.4]
  assign _T_10181 = offsetQ_10 < 4'h5; // @[LoadQueue.scala 132:33:@10512.4]
  assign _T_10184 = _T_10181 & _T_6217; // @[LoadQueue.scala 132:41:@10514.4]
  assign _T_10186 = _T_10184 == 1'h0; // @[LoadQueue.scala 132:9:@10515.4]
  assign storesToCheck_10_5 = _T_2536 ? _T_10179 : _T_10186; // @[LoadQueue.scala 131:10:@10516.4]
  assign _T_10192 = 4'h6 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10519.4]
  assign _T_10193 = _T_6225 & _T_10192; // @[LoadQueue.scala 131:72:@10520.4]
  assign _T_10195 = offsetQ_10 < 4'h6; // @[LoadQueue.scala 132:33:@10521.4]
  assign _T_10198 = _T_10195 & _T_6234; // @[LoadQueue.scala 132:41:@10523.4]
  assign _T_10200 = _T_10198 == 1'h0; // @[LoadQueue.scala 132:9:@10524.4]
  assign storesToCheck_10_6 = _T_2536 ? _T_10193 : _T_10200; // @[LoadQueue.scala 131:10:@10525.4]
  assign _T_10206 = 4'h7 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10528.4]
  assign _T_10207 = _T_6242 & _T_10206; // @[LoadQueue.scala 131:72:@10529.4]
  assign _T_10209 = offsetQ_10 < 4'h7; // @[LoadQueue.scala 132:33:@10530.4]
  assign _T_10212 = _T_10209 & _T_6251; // @[LoadQueue.scala 132:41:@10532.4]
  assign _T_10214 = _T_10212 == 1'h0; // @[LoadQueue.scala 132:9:@10533.4]
  assign storesToCheck_10_7 = _T_2536 ? _T_10207 : _T_10214; // @[LoadQueue.scala 131:10:@10534.4]
  assign _T_10220 = 4'h8 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10537.4]
  assign _T_10221 = _T_6259 & _T_10220; // @[LoadQueue.scala 131:72:@10538.4]
  assign _T_10223 = offsetQ_10 < 4'h8; // @[LoadQueue.scala 132:33:@10539.4]
  assign _T_10226 = _T_10223 & _T_6268; // @[LoadQueue.scala 132:41:@10541.4]
  assign _T_10228 = _T_10226 == 1'h0; // @[LoadQueue.scala 132:9:@10542.4]
  assign storesToCheck_10_8 = _T_2536 ? _T_10221 : _T_10228; // @[LoadQueue.scala 131:10:@10543.4]
  assign _T_10234 = 4'h9 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10546.4]
  assign _T_10235 = _T_6276 & _T_10234; // @[LoadQueue.scala 131:72:@10547.4]
  assign _T_10237 = offsetQ_10 < 4'h9; // @[LoadQueue.scala 132:33:@10548.4]
  assign _T_10240 = _T_10237 & _T_6285; // @[LoadQueue.scala 132:41:@10550.4]
  assign _T_10242 = _T_10240 == 1'h0; // @[LoadQueue.scala 132:9:@10551.4]
  assign storesToCheck_10_9 = _T_2536 ? _T_10235 : _T_10242; // @[LoadQueue.scala 131:10:@10552.4]
  assign _T_10248 = 4'ha <= offsetQ_10; // @[LoadQueue.scala 131:81:@10555.4]
  assign _T_10249 = _T_6293 & _T_10248; // @[LoadQueue.scala 131:72:@10556.4]
  assign _T_10251 = offsetQ_10 < 4'ha; // @[LoadQueue.scala 132:33:@10557.4]
  assign _T_10254 = _T_10251 & _T_6302; // @[LoadQueue.scala 132:41:@10559.4]
  assign _T_10256 = _T_10254 == 1'h0; // @[LoadQueue.scala 132:9:@10560.4]
  assign storesToCheck_10_10 = _T_2536 ? _T_10249 : _T_10256; // @[LoadQueue.scala 131:10:@10561.4]
  assign _T_10262 = 4'hb <= offsetQ_10; // @[LoadQueue.scala 131:81:@10564.4]
  assign _T_10263 = _T_6310 & _T_10262; // @[LoadQueue.scala 131:72:@10565.4]
  assign _T_10265 = offsetQ_10 < 4'hb; // @[LoadQueue.scala 132:33:@10566.4]
  assign _T_10268 = _T_10265 & _T_6319; // @[LoadQueue.scala 132:41:@10568.4]
  assign _T_10270 = _T_10268 == 1'h0; // @[LoadQueue.scala 132:9:@10569.4]
  assign storesToCheck_10_11 = _T_2536 ? _T_10263 : _T_10270; // @[LoadQueue.scala 131:10:@10570.4]
  assign _T_10276 = 4'hc <= offsetQ_10; // @[LoadQueue.scala 131:81:@10573.4]
  assign _T_10277 = _T_6327 & _T_10276; // @[LoadQueue.scala 131:72:@10574.4]
  assign _T_10279 = offsetQ_10 < 4'hc; // @[LoadQueue.scala 132:33:@10575.4]
  assign _T_10282 = _T_10279 & _T_6336; // @[LoadQueue.scala 132:41:@10577.4]
  assign _T_10284 = _T_10282 == 1'h0; // @[LoadQueue.scala 132:9:@10578.4]
  assign storesToCheck_10_12 = _T_2536 ? _T_10277 : _T_10284; // @[LoadQueue.scala 131:10:@10579.4]
  assign _T_10290 = 4'hd <= offsetQ_10; // @[LoadQueue.scala 131:81:@10582.4]
  assign _T_10291 = _T_6344 & _T_10290; // @[LoadQueue.scala 131:72:@10583.4]
  assign _T_10293 = offsetQ_10 < 4'hd; // @[LoadQueue.scala 132:33:@10584.4]
  assign _T_10296 = _T_10293 & _T_6353; // @[LoadQueue.scala 132:41:@10586.4]
  assign _T_10298 = _T_10296 == 1'h0; // @[LoadQueue.scala 132:9:@10587.4]
  assign storesToCheck_10_13 = _T_2536 ? _T_10291 : _T_10298; // @[LoadQueue.scala 131:10:@10588.4]
  assign _T_10304 = 4'he <= offsetQ_10; // @[LoadQueue.scala 131:81:@10591.4]
  assign _T_10305 = _T_6361 & _T_10304; // @[LoadQueue.scala 131:72:@10592.4]
  assign _T_10307 = offsetQ_10 < 4'he; // @[LoadQueue.scala 132:33:@10593.4]
  assign _T_10310 = _T_10307 & _T_6370; // @[LoadQueue.scala 132:41:@10595.4]
  assign _T_10312 = _T_10310 == 1'h0; // @[LoadQueue.scala 132:9:@10596.4]
  assign storesToCheck_10_14 = _T_2536 ? _T_10305 : _T_10312; // @[LoadQueue.scala 131:10:@10597.4]
  assign _T_10318 = 4'hf <= offsetQ_10; // @[LoadQueue.scala 131:81:@10600.4]
  assign storesToCheck_10_15 = _T_2536 ? _T_10318 : 1'h1; // @[LoadQueue.scala 131:10:@10606.4]
  assign storesToCheck_11_0 = _T_2566 ? _T_6123 : 1'h1; // @[LoadQueue.scala 131:10:@10648.4]
  assign _T_10368 = 4'h1 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10651.4]
  assign _T_10369 = _T_6140 & _T_10368; // @[LoadQueue.scala 131:72:@10652.4]
  assign _T_10371 = offsetQ_11 < 4'h1; // @[LoadQueue.scala 132:33:@10653.4]
  assign _T_10374 = _T_10371 & _T_6149; // @[LoadQueue.scala 132:41:@10655.4]
  assign _T_10376 = _T_10374 == 1'h0; // @[LoadQueue.scala 132:9:@10656.4]
  assign storesToCheck_11_1 = _T_2566 ? _T_10369 : _T_10376; // @[LoadQueue.scala 131:10:@10657.4]
  assign _T_10382 = 4'h2 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10660.4]
  assign _T_10383 = _T_6157 & _T_10382; // @[LoadQueue.scala 131:72:@10661.4]
  assign _T_10385 = offsetQ_11 < 4'h2; // @[LoadQueue.scala 132:33:@10662.4]
  assign _T_10388 = _T_10385 & _T_6166; // @[LoadQueue.scala 132:41:@10664.4]
  assign _T_10390 = _T_10388 == 1'h0; // @[LoadQueue.scala 132:9:@10665.4]
  assign storesToCheck_11_2 = _T_2566 ? _T_10383 : _T_10390; // @[LoadQueue.scala 131:10:@10666.4]
  assign _T_10396 = 4'h3 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10669.4]
  assign _T_10397 = _T_6174 & _T_10396; // @[LoadQueue.scala 131:72:@10670.4]
  assign _T_10399 = offsetQ_11 < 4'h3; // @[LoadQueue.scala 132:33:@10671.4]
  assign _T_10402 = _T_10399 & _T_6183; // @[LoadQueue.scala 132:41:@10673.4]
  assign _T_10404 = _T_10402 == 1'h0; // @[LoadQueue.scala 132:9:@10674.4]
  assign storesToCheck_11_3 = _T_2566 ? _T_10397 : _T_10404; // @[LoadQueue.scala 131:10:@10675.4]
  assign _T_10410 = 4'h4 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10678.4]
  assign _T_10411 = _T_6191 & _T_10410; // @[LoadQueue.scala 131:72:@10679.4]
  assign _T_10413 = offsetQ_11 < 4'h4; // @[LoadQueue.scala 132:33:@10680.4]
  assign _T_10416 = _T_10413 & _T_6200; // @[LoadQueue.scala 132:41:@10682.4]
  assign _T_10418 = _T_10416 == 1'h0; // @[LoadQueue.scala 132:9:@10683.4]
  assign storesToCheck_11_4 = _T_2566 ? _T_10411 : _T_10418; // @[LoadQueue.scala 131:10:@10684.4]
  assign _T_10424 = 4'h5 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10687.4]
  assign _T_10425 = _T_6208 & _T_10424; // @[LoadQueue.scala 131:72:@10688.4]
  assign _T_10427 = offsetQ_11 < 4'h5; // @[LoadQueue.scala 132:33:@10689.4]
  assign _T_10430 = _T_10427 & _T_6217; // @[LoadQueue.scala 132:41:@10691.4]
  assign _T_10432 = _T_10430 == 1'h0; // @[LoadQueue.scala 132:9:@10692.4]
  assign storesToCheck_11_5 = _T_2566 ? _T_10425 : _T_10432; // @[LoadQueue.scala 131:10:@10693.4]
  assign _T_10438 = 4'h6 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10696.4]
  assign _T_10439 = _T_6225 & _T_10438; // @[LoadQueue.scala 131:72:@10697.4]
  assign _T_10441 = offsetQ_11 < 4'h6; // @[LoadQueue.scala 132:33:@10698.4]
  assign _T_10444 = _T_10441 & _T_6234; // @[LoadQueue.scala 132:41:@10700.4]
  assign _T_10446 = _T_10444 == 1'h0; // @[LoadQueue.scala 132:9:@10701.4]
  assign storesToCheck_11_6 = _T_2566 ? _T_10439 : _T_10446; // @[LoadQueue.scala 131:10:@10702.4]
  assign _T_10452 = 4'h7 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10705.4]
  assign _T_10453 = _T_6242 & _T_10452; // @[LoadQueue.scala 131:72:@10706.4]
  assign _T_10455 = offsetQ_11 < 4'h7; // @[LoadQueue.scala 132:33:@10707.4]
  assign _T_10458 = _T_10455 & _T_6251; // @[LoadQueue.scala 132:41:@10709.4]
  assign _T_10460 = _T_10458 == 1'h0; // @[LoadQueue.scala 132:9:@10710.4]
  assign storesToCheck_11_7 = _T_2566 ? _T_10453 : _T_10460; // @[LoadQueue.scala 131:10:@10711.4]
  assign _T_10466 = 4'h8 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10714.4]
  assign _T_10467 = _T_6259 & _T_10466; // @[LoadQueue.scala 131:72:@10715.4]
  assign _T_10469 = offsetQ_11 < 4'h8; // @[LoadQueue.scala 132:33:@10716.4]
  assign _T_10472 = _T_10469 & _T_6268; // @[LoadQueue.scala 132:41:@10718.4]
  assign _T_10474 = _T_10472 == 1'h0; // @[LoadQueue.scala 132:9:@10719.4]
  assign storesToCheck_11_8 = _T_2566 ? _T_10467 : _T_10474; // @[LoadQueue.scala 131:10:@10720.4]
  assign _T_10480 = 4'h9 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10723.4]
  assign _T_10481 = _T_6276 & _T_10480; // @[LoadQueue.scala 131:72:@10724.4]
  assign _T_10483 = offsetQ_11 < 4'h9; // @[LoadQueue.scala 132:33:@10725.4]
  assign _T_10486 = _T_10483 & _T_6285; // @[LoadQueue.scala 132:41:@10727.4]
  assign _T_10488 = _T_10486 == 1'h0; // @[LoadQueue.scala 132:9:@10728.4]
  assign storesToCheck_11_9 = _T_2566 ? _T_10481 : _T_10488; // @[LoadQueue.scala 131:10:@10729.4]
  assign _T_10494 = 4'ha <= offsetQ_11; // @[LoadQueue.scala 131:81:@10732.4]
  assign _T_10495 = _T_6293 & _T_10494; // @[LoadQueue.scala 131:72:@10733.4]
  assign _T_10497 = offsetQ_11 < 4'ha; // @[LoadQueue.scala 132:33:@10734.4]
  assign _T_10500 = _T_10497 & _T_6302; // @[LoadQueue.scala 132:41:@10736.4]
  assign _T_10502 = _T_10500 == 1'h0; // @[LoadQueue.scala 132:9:@10737.4]
  assign storesToCheck_11_10 = _T_2566 ? _T_10495 : _T_10502; // @[LoadQueue.scala 131:10:@10738.4]
  assign _T_10508 = 4'hb <= offsetQ_11; // @[LoadQueue.scala 131:81:@10741.4]
  assign _T_10509 = _T_6310 & _T_10508; // @[LoadQueue.scala 131:72:@10742.4]
  assign _T_10511 = offsetQ_11 < 4'hb; // @[LoadQueue.scala 132:33:@10743.4]
  assign _T_10514 = _T_10511 & _T_6319; // @[LoadQueue.scala 132:41:@10745.4]
  assign _T_10516 = _T_10514 == 1'h0; // @[LoadQueue.scala 132:9:@10746.4]
  assign storesToCheck_11_11 = _T_2566 ? _T_10509 : _T_10516; // @[LoadQueue.scala 131:10:@10747.4]
  assign _T_10522 = 4'hc <= offsetQ_11; // @[LoadQueue.scala 131:81:@10750.4]
  assign _T_10523 = _T_6327 & _T_10522; // @[LoadQueue.scala 131:72:@10751.4]
  assign _T_10525 = offsetQ_11 < 4'hc; // @[LoadQueue.scala 132:33:@10752.4]
  assign _T_10528 = _T_10525 & _T_6336; // @[LoadQueue.scala 132:41:@10754.4]
  assign _T_10530 = _T_10528 == 1'h0; // @[LoadQueue.scala 132:9:@10755.4]
  assign storesToCheck_11_12 = _T_2566 ? _T_10523 : _T_10530; // @[LoadQueue.scala 131:10:@10756.4]
  assign _T_10536 = 4'hd <= offsetQ_11; // @[LoadQueue.scala 131:81:@10759.4]
  assign _T_10537 = _T_6344 & _T_10536; // @[LoadQueue.scala 131:72:@10760.4]
  assign _T_10539 = offsetQ_11 < 4'hd; // @[LoadQueue.scala 132:33:@10761.4]
  assign _T_10542 = _T_10539 & _T_6353; // @[LoadQueue.scala 132:41:@10763.4]
  assign _T_10544 = _T_10542 == 1'h0; // @[LoadQueue.scala 132:9:@10764.4]
  assign storesToCheck_11_13 = _T_2566 ? _T_10537 : _T_10544; // @[LoadQueue.scala 131:10:@10765.4]
  assign _T_10550 = 4'he <= offsetQ_11; // @[LoadQueue.scala 131:81:@10768.4]
  assign _T_10551 = _T_6361 & _T_10550; // @[LoadQueue.scala 131:72:@10769.4]
  assign _T_10553 = offsetQ_11 < 4'he; // @[LoadQueue.scala 132:33:@10770.4]
  assign _T_10556 = _T_10553 & _T_6370; // @[LoadQueue.scala 132:41:@10772.4]
  assign _T_10558 = _T_10556 == 1'h0; // @[LoadQueue.scala 132:9:@10773.4]
  assign storesToCheck_11_14 = _T_2566 ? _T_10551 : _T_10558; // @[LoadQueue.scala 131:10:@10774.4]
  assign _T_10564 = 4'hf <= offsetQ_11; // @[LoadQueue.scala 131:81:@10777.4]
  assign storesToCheck_11_15 = _T_2566 ? _T_10564 : 1'h1; // @[LoadQueue.scala 131:10:@10783.4]
  assign storesToCheck_12_0 = _T_2596 ? _T_6123 : 1'h1; // @[LoadQueue.scala 131:10:@10825.4]
  assign _T_10614 = 4'h1 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10828.4]
  assign _T_10615 = _T_6140 & _T_10614; // @[LoadQueue.scala 131:72:@10829.4]
  assign _T_10617 = offsetQ_12 < 4'h1; // @[LoadQueue.scala 132:33:@10830.4]
  assign _T_10620 = _T_10617 & _T_6149; // @[LoadQueue.scala 132:41:@10832.4]
  assign _T_10622 = _T_10620 == 1'h0; // @[LoadQueue.scala 132:9:@10833.4]
  assign storesToCheck_12_1 = _T_2596 ? _T_10615 : _T_10622; // @[LoadQueue.scala 131:10:@10834.4]
  assign _T_10628 = 4'h2 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10837.4]
  assign _T_10629 = _T_6157 & _T_10628; // @[LoadQueue.scala 131:72:@10838.4]
  assign _T_10631 = offsetQ_12 < 4'h2; // @[LoadQueue.scala 132:33:@10839.4]
  assign _T_10634 = _T_10631 & _T_6166; // @[LoadQueue.scala 132:41:@10841.4]
  assign _T_10636 = _T_10634 == 1'h0; // @[LoadQueue.scala 132:9:@10842.4]
  assign storesToCheck_12_2 = _T_2596 ? _T_10629 : _T_10636; // @[LoadQueue.scala 131:10:@10843.4]
  assign _T_10642 = 4'h3 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10846.4]
  assign _T_10643 = _T_6174 & _T_10642; // @[LoadQueue.scala 131:72:@10847.4]
  assign _T_10645 = offsetQ_12 < 4'h3; // @[LoadQueue.scala 132:33:@10848.4]
  assign _T_10648 = _T_10645 & _T_6183; // @[LoadQueue.scala 132:41:@10850.4]
  assign _T_10650 = _T_10648 == 1'h0; // @[LoadQueue.scala 132:9:@10851.4]
  assign storesToCheck_12_3 = _T_2596 ? _T_10643 : _T_10650; // @[LoadQueue.scala 131:10:@10852.4]
  assign _T_10656 = 4'h4 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10855.4]
  assign _T_10657 = _T_6191 & _T_10656; // @[LoadQueue.scala 131:72:@10856.4]
  assign _T_10659 = offsetQ_12 < 4'h4; // @[LoadQueue.scala 132:33:@10857.4]
  assign _T_10662 = _T_10659 & _T_6200; // @[LoadQueue.scala 132:41:@10859.4]
  assign _T_10664 = _T_10662 == 1'h0; // @[LoadQueue.scala 132:9:@10860.4]
  assign storesToCheck_12_4 = _T_2596 ? _T_10657 : _T_10664; // @[LoadQueue.scala 131:10:@10861.4]
  assign _T_10670 = 4'h5 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10864.4]
  assign _T_10671 = _T_6208 & _T_10670; // @[LoadQueue.scala 131:72:@10865.4]
  assign _T_10673 = offsetQ_12 < 4'h5; // @[LoadQueue.scala 132:33:@10866.4]
  assign _T_10676 = _T_10673 & _T_6217; // @[LoadQueue.scala 132:41:@10868.4]
  assign _T_10678 = _T_10676 == 1'h0; // @[LoadQueue.scala 132:9:@10869.4]
  assign storesToCheck_12_5 = _T_2596 ? _T_10671 : _T_10678; // @[LoadQueue.scala 131:10:@10870.4]
  assign _T_10684 = 4'h6 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10873.4]
  assign _T_10685 = _T_6225 & _T_10684; // @[LoadQueue.scala 131:72:@10874.4]
  assign _T_10687 = offsetQ_12 < 4'h6; // @[LoadQueue.scala 132:33:@10875.4]
  assign _T_10690 = _T_10687 & _T_6234; // @[LoadQueue.scala 132:41:@10877.4]
  assign _T_10692 = _T_10690 == 1'h0; // @[LoadQueue.scala 132:9:@10878.4]
  assign storesToCheck_12_6 = _T_2596 ? _T_10685 : _T_10692; // @[LoadQueue.scala 131:10:@10879.4]
  assign _T_10698 = 4'h7 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10882.4]
  assign _T_10699 = _T_6242 & _T_10698; // @[LoadQueue.scala 131:72:@10883.4]
  assign _T_10701 = offsetQ_12 < 4'h7; // @[LoadQueue.scala 132:33:@10884.4]
  assign _T_10704 = _T_10701 & _T_6251; // @[LoadQueue.scala 132:41:@10886.4]
  assign _T_10706 = _T_10704 == 1'h0; // @[LoadQueue.scala 132:9:@10887.4]
  assign storesToCheck_12_7 = _T_2596 ? _T_10699 : _T_10706; // @[LoadQueue.scala 131:10:@10888.4]
  assign _T_10712 = 4'h8 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10891.4]
  assign _T_10713 = _T_6259 & _T_10712; // @[LoadQueue.scala 131:72:@10892.4]
  assign _T_10715 = offsetQ_12 < 4'h8; // @[LoadQueue.scala 132:33:@10893.4]
  assign _T_10718 = _T_10715 & _T_6268; // @[LoadQueue.scala 132:41:@10895.4]
  assign _T_10720 = _T_10718 == 1'h0; // @[LoadQueue.scala 132:9:@10896.4]
  assign storesToCheck_12_8 = _T_2596 ? _T_10713 : _T_10720; // @[LoadQueue.scala 131:10:@10897.4]
  assign _T_10726 = 4'h9 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10900.4]
  assign _T_10727 = _T_6276 & _T_10726; // @[LoadQueue.scala 131:72:@10901.4]
  assign _T_10729 = offsetQ_12 < 4'h9; // @[LoadQueue.scala 132:33:@10902.4]
  assign _T_10732 = _T_10729 & _T_6285; // @[LoadQueue.scala 132:41:@10904.4]
  assign _T_10734 = _T_10732 == 1'h0; // @[LoadQueue.scala 132:9:@10905.4]
  assign storesToCheck_12_9 = _T_2596 ? _T_10727 : _T_10734; // @[LoadQueue.scala 131:10:@10906.4]
  assign _T_10740 = 4'ha <= offsetQ_12; // @[LoadQueue.scala 131:81:@10909.4]
  assign _T_10741 = _T_6293 & _T_10740; // @[LoadQueue.scala 131:72:@10910.4]
  assign _T_10743 = offsetQ_12 < 4'ha; // @[LoadQueue.scala 132:33:@10911.4]
  assign _T_10746 = _T_10743 & _T_6302; // @[LoadQueue.scala 132:41:@10913.4]
  assign _T_10748 = _T_10746 == 1'h0; // @[LoadQueue.scala 132:9:@10914.4]
  assign storesToCheck_12_10 = _T_2596 ? _T_10741 : _T_10748; // @[LoadQueue.scala 131:10:@10915.4]
  assign _T_10754 = 4'hb <= offsetQ_12; // @[LoadQueue.scala 131:81:@10918.4]
  assign _T_10755 = _T_6310 & _T_10754; // @[LoadQueue.scala 131:72:@10919.4]
  assign _T_10757 = offsetQ_12 < 4'hb; // @[LoadQueue.scala 132:33:@10920.4]
  assign _T_10760 = _T_10757 & _T_6319; // @[LoadQueue.scala 132:41:@10922.4]
  assign _T_10762 = _T_10760 == 1'h0; // @[LoadQueue.scala 132:9:@10923.4]
  assign storesToCheck_12_11 = _T_2596 ? _T_10755 : _T_10762; // @[LoadQueue.scala 131:10:@10924.4]
  assign _T_10768 = 4'hc <= offsetQ_12; // @[LoadQueue.scala 131:81:@10927.4]
  assign _T_10769 = _T_6327 & _T_10768; // @[LoadQueue.scala 131:72:@10928.4]
  assign _T_10771 = offsetQ_12 < 4'hc; // @[LoadQueue.scala 132:33:@10929.4]
  assign _T_10774 = _T_10771 & _T_6336; // @[LoadQueue.scala 132:41:@10931.4]
  assign _T_10776 = _T_10774 == 1'h0; // @[LoadQueue.scala 132:9:@10932.4]
  assign storesToCheck_12_12 = _T_2596 ? _T_10769 : _T_10776; // @[LoadQueue.scala 131:10:@10933.4]
  assign _T_10782 = 4'hd <= offsetQ_12; // @[LoadQueue.scala 131:81:@10936.4]
  assign _T_10783 = _T_6344 & _T_10782; // @[LoadQueue.scala 131:72:@10937.4]
  assign _T_10785 = offsetQ_12 < 4'hd; // @[LoadQueue.scala 132:33:@10938.4]
  assign _T_10788 = _T_10785 & _T_6353; // @[LoadQueue.scala 132:41:@10940.4]
  assign _T_10790 = _T_10788 == 1'h0; // @[LoadQueue.scala 132:9:@10941.4]
  assign storesToCheck_12_13 = _T_2596 ? _T_10783 : _T_10790; // @[LoadQueue.scala 131:10:@10942.4]
  assign _T_10796 = 4'he <= offsetQ_12; // @[LoadQueue.scala 131:81:@10945.4]
  assign _T_10797 = _T_6361 & _T_10796; // @[LoadQueue.scala 131:72:@10946.4]
  assign _T_10799 = offsetQ_12 < 4'he; // @[LoadQueue.scala 132:33:@10947.4]
  assign _T_10802 = _T_10799 & _T_6370; // @[LoadQueue.scala 132:41:@10949.4]
  assign _T_10804 = _T_10802 == 1'h0; // @[LoadQueue.scala 132:9:@10950.4]
  assign storesToCheck_12_14 = _T_2596 ? _T_10797 : _T_10804; // @[LoadQueue.scala 131:10:@10951.4]
  assign _T_10810 = 4'hf <= offsetQ_12; // @[LoadQueue.scala 131:81:@10954.4]
  assign storesToCheck_12_15 = _T_2596 ? _T_10810 : 1'h1; // @[LoadQueue.scala 131:10:@10960.4]
  assign storesToCheck_13_0 = _T_2626 ? _T_6123 : 1'h1; // @[LoadQueue.scala 131:10:@11002.4]
  assign _T_10860 = 4'h1 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11005.4]
  assign _T_10861 = _T_6140 & _T_10860; // @[LoadQueue.scala 131:72:@11006.4]
  assign _T_10863 = offsetQ_13 < 4'h1; // @[LoadQueue.scala 132:33:@11007.4]
  assign _T_10866 = _T_10863 & _T_6149; // @[LoadQueue.scala 132:41:@11009.4]
  assign _T_10868 = _T_10866 == 1'h0; // @[LoadQueue.scala 132:9:@11010.4]
  assign storesToCheck_13_1 = _T_2626 ? _T_10861 : _T_10868; // @[LoadQueue.scala 131:10:@11011.4]
  assign _T_10874 = 4'h2 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11014.4]
  assign _T_10875 = _T_6157 & _T_10874; // @[LoadQueue.scala 131:72:@11015.4]
  assign _T_10877 = offsetQ_13 < 4'h2; // @[LoadQueue.scala 132:33:@11016.4]
  assign _T_10880 = _T_10877 & _T_6166; // @[LoadQueue.scala 132:41:@11018.4]
  assign _T_10882 = _T_10880 == 1'h0; // @[LoadQueue.scala 132:9:@11019.4]
  assign storesToCheck_13_2 = _T_2626 ? _T_10875 : _T_10882; // @[LoadQueue.scala 131:10:@11020.4]
  assign _T_10888 = 4'h3 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11023.4]
  assign _T_10889 = _T_6174 & _T_10888; // @[LoadQueue.scala 131:72:@11024.4]
  assign _T_10891 = offsetQ_13 < 4'h3; // @[LoadQueue.scala 132:33:@11025.4]
  assign _T_10894 = _T_10891 & _T_6183; // @[LoadQueue.scala 132:41:@11027.4]
  assign _T_10896 = _T_10894 == 1'h0; // @[LoadQueue.scala 132:9:@11028.4]
  assign storesToCheck_13_3 = _T_2626 ? _T_10889 : _T_10896; // @[LoadQueue.scala 131:10:@11029.4]
  assign _T_10902 = 4'h4 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11032.4]
  assign _T_10903 = _T_6191 & _T_10902; // @[LoadQueue.scala 131:72:@11033.4]
  assign _T_10905 = offsetQ_13 < 4'h4; // @[LoadQueue.scala 132:33:@11034.4]
  assign _T_10908 = _T_10905 & _T_6200; // @[LoadQueue.scala 132:41:@11036.4]
  assign _T_10910 = _T_10908 == 1'h0; // @[LoadQueue.scala 132:9:@11037.4]
  assign storesToCheck_13_4 = _T_2626 ? _T_10903 : _T_10910; // @[LoadQueue.scala 131:10:@11038.4]
  assign _T_10916 = 4'h5 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11041.4]
  assign _T_10917 = _T_6208 & _T_10916; // @[LoadQueue.scala 131:72:@11042.4]
  assign _T_10919 = offsetQ_13 < 4'h5; // @[LoadQueue.scala 132:33:@11043.4]
  assign _T_10922 = _T_10919 & _T_6217; // @[LoadQueue.scala 132:41:@11045.4]
  assign _T_10924 = _T_10922 == 1'h0; // @[LoadQueue.scala 132:9:@11046.4]
  assign storesToCheck_13_5 = _T_2626 ? _T_10917 : _T_10924; // @[LoadQueue.scala 131:10:@11047.4]
  assign _T_10930 = 4'h6 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11050.4]
  assign _T_10931 = _T_6225 & _T_10930; // @[LoadQueue.scala 131:72:@11051.4]
  assign _T_10933 = offsetQ_13 < 4'h6; // @[LoadQueue.scala 132:33:@11052.4]
  assign _T_10936 = _T_10933 & _T_6234; // @[LoadQueue.scala 132:41:@11054.4]
  assign _T_10938 = _T_10936 == 1'h0; // @[LoadQueue.scala 132:9:@11055.4]
  assign storesToCheck_13_6 = _T_2626 ? _T_10931 : _T_10938; // @[LoadQueue.scala 131:10:@11056.4]
  assign _T_10944 = 4'h7 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11059.4]
  assign _T_10945 = _T_6242 & _T_10944; // @[LoadQueue.scala 131:72:@11060.4]
  assign _T_10947 = offsetQ_13 < 4'h7; // @[LoadQueue.scala 132:33:@11061.4]
  assign _T_10950 = _T_10947 & _T_6251; // @[LoadQueue.scala 132:41:@11063.4]
  assign _T_10952 = _T_10950 == 1'h0; // @[LoadQueue.scala 132:9:@11064.4]
  assign storesToCheck_13_7 = _T_2626 ? _T_10945 : _T_10952; // @[LoadQueue.scala 131:10:@11065.4]
  assign _T_10958 = 4'h8 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11068.4]
  assign _T_10959 = _T_6259 & _T_10958; // @[LoadQueue.scala 131:72:@11069.4]
  assign _T_10961 = offsetQ_13 < 4'h8; // @[LoadQueue.scala 132:33:@11070.4]
  assign _T_10964 = _T_10961 & _T_6268; // @[LoadQueue.scala 132:41:@11072.4]
  assign _T_10966 = _T_10964 == 1'h0; // @[LoadQueue.scala 132:9:@11073.4]
  assign storesToCheck_13_8 = _T_2626 ? _T_10959 : _T_10966; // @[LoadQueue.scala 131:10:@11074.4]
  assign _T_10972 = 4'h9 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11077.4]
  assign _T_10973 = _T_6276 & _T_10972; // @[LoadQueue.scala 131:72:@11078.4]
  assign _T_10975 = offsetQ_13 < 4'h9; // @[LoadQueue.scala 132:33:@11079.4]
  assign _T_10978 = _T_10975 & _T_6285; // @[LoadQueue.scala 132:41:@11081.4]
  assign _T_10980 = _T_10978 == 1'h0; // @[LoadQueue.scala 132:9:@11082.4]
  assign storesToCheck_13_9 = _T_2626 ? _T_10973 : _T_10980; // @[LoadQueue.scala 131:10:@11083.4]
  assign _T_10986 = 4'ha <= offsetQ_13; // @[LoadQueue.scala 131:81:@11086.4]
  assign _T_10987 = _T_6293 & _T_10986; // @[LoadQueue.scala 131:72:@11087.4]
  assign _T_10989 = offsetQ_13 < 4'ha; // @[LoadQueue.scala 132:33:@11088.4]
  assign _T_10992 = _T_10989 & _T_6302; // @[LoadQueue.scala 132:41:@11090.4]
  assign _T_10994 = _T_10992 == 1'h0; // @[LoadQueue.scala 132:9:@11091.4]
  assign storesToCheck_13_10 = _T_2626 ? _T_10987 : _T_10994; // @[LoadQueue.scala 131:10:@11092.4]
  assign _T_11000 = 4'hb <= offsetQ_13; // @[LoadQueue.scala 131:81:@11095.4]
  assign _T_11001 = _T_6310 & _T_11000; // @[LoadQueue.scala 131:72:@11096.4]
  assign _T_11003 = offsetQ_13 < 4'hb; // @[LoadQueue.scala 132:33:@11097.4]
  assign _T_11006 = _T_11003 & _T_6319; // @[LoadQueue.scala 132:41:@11099.4]
  assign _T_11008 = _T_11006 == 1'h0; // @[LoadQueue.scala 132:9:@11100.4]
  assign storesToCheck_13_11 = _T_2626 ? _T_11001 : _T_11008; // @[LoadQueue.scala 131:10:@11101.4]
  assign _T_11014 = 4'hc <= offsetQ_13; // @[LoadQueue.scala 131:81:@11104.4]
  assign _T_11015 = _T_6327 & _T_11014; // @[LoadQueue.scala 131:72:@11105.4]
  assign _T_11017 = offsetQ_13 < 4'hc; // @[LoadQueue.scala 132:33:@11106.4]
  assign _T_11020 = _T_11017 & _T_6336; // @[LoadQueue.scala 132:41:@11108.4]
  assign _T_11022 = _T_11020 == 1'h0; // @[LoadQueue.scala 132:9:@11109.4]
  assign storesToCheck_13_12 = _T_2626 ? _T_11015 : _T_11022; // @[LoadQueue.scala 131:10:@11110.4]
  assign _T_11028 = 4'hd <= offsetQ_13; // @[LoadQueue.scala 131:81:@11113.4]
  assign _T_11029 = _T_6344 & _T_11028; // @[LoadQueue.scala 131:72:@11114.4]
  assign _T_11031 = offsetQ_13 < 4'hd; // @[LoadQueue.scala 132:33:@11115.4]
  assign _T_11034 = _T_11031 & _T_6353; // @[LoadQueue.scala 132:41:@11117.4]
  assign _T_11036 = _T_11034 == 1'h0; // @[LoadQueue.scala 132:9:@11118.4]
  assign storesToCheck_13_13 = _T_2626 ? _T_11029 : _T_11036; // @[LoadQueue.scala 131:10:@11119.4]
  assign _T_11042 = 4'he <= offsetQ_13; // @[LoadQueue.scala 131:81:@11122.4]
  assign _T_11043 = _T_6361 & _T_11042; // @[LoadQueue.scala 131:72:@11123.4]
  assign _T_11045 = offsetQ_13 < 4'he; // @[LoadQueue.scala 132:33:@11124.4]
  assign _T_11048 = _T_11045 & _T_6370; // @[LoadQueue.scala 132:41:@11126.4]
  assign _T_11050 = _T_11048 == 1'h0; // @[LoadQueue.scala 132:9:@11127.4]
  assign storesToCheck_13_14 = _T_2626 ? _T_11043 : _T_11050; // @[LoadQueue.scala 131:10:@11128.4]
  assign _T_11056 = 4'hf <= offsetQ_13; // @[LoadQueue.scala 131:81:@11131.4]
  assign storesToCheck_13_15 = _T_2626 ? _T_11056 : 1'h1; // @[LoadQueue.scala 131:10:@11137.4]
  assign storesToCheck_14_0 = _T_2656 ? _T_6123 : 1'h1; // @[LoadQueue.scala 131:10:@11179.4]
  assign _T_11106 = 4'h1 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11182.4]
  assign _T_11107 = _T_6140 & _T_11106; // @[LoadQueue.scala 131:72:@11183.4]
  assign _T_11109 = offsetQ_14 < 4'h1; // @[LoadQueue.scala 132:33:@11184.4]
  assign _T_11112 = _T_11109 & _T_6149; // @[LoadQueue.scala 132:41:@11186.4]
  assign _T_11114 = _T_11112 == 1'h0; // @[LoadQueue.scala 132:9:@11187.4]
  assign storesToCheck_14_1 = _T_2656 ? _T_11107 : _T_11114; // @[LoadQueue.scala 131:10:@11188.4]
  assign _T_11120 = 4'h2 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11191.4]
  assign _T_11121 = _T_6157 & _T_11120; // @[LoadQueue.scala 131:72:@11192.4]
  assign _T_11123 = offsetQ_14 < 4'h2; // @[LoadQueue.scala 132:33:@11193.4]
  assign _T_11126 = _T_11123 & _T_6166; // @[LoadQueue.scala 132:41:@11195.4]
  assign _T_11128 = _T_11126 == 1'h0; // @[LoadQueue.scala 132:9:@11196.4]
  assign storesToCheck_14_2 = _T_2656 ? _T_11121 : _T_11128; // @[LoadQueue.scala 131:10:@11197.4]
  assign _T_11134 = 4'h3 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11200.4]
  assign _T_11135 = _T_6174 & _T_11134; // @[LoadQueue.scala 131:72:@11201.4]
  assign _T_11137 = offsetQ_14 < 4'h3; // @[LoadQueue.scala 132:33:@11202.4]
  assign _T_11140 = _T_11137 & _T_6183; // @[LoadQueue.scala 132:41:@11204.4]
  assign _T_11142 = _T_11140 == 1'h0; // @[LoadQueue.scala 132:9:@11205.4]
  assign storesToCheck_14_3 = _T_2656 ? _T_11135 : _T_11142; // @[LoadQueue.scala 131:10:@11206.4]
  assign _T_11148 = 4'h4 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11209.4]
  assign _T_11149 = _T_6191 & _T_11148; // @[LoadQueue.scala 131:72:@11210.4]
  assign _T_11151 = offsetQ_14 < 4'h4; // @[LoadQueue.scala 132:33:@11211.4]
  assign _T_11154 = _T_11151 & _T_6200; // @[LoadQueue.scala 132:41:@11213.4]
  assign _T_11156 = _T_11154 == 1'h0; // @[LoadQueue.scala 132:9:@11214.4]
  assign storesToCheck_14_4 = _T_2656 ? _T_11149 : _T_11156; // @[LoadQueue.scala 131:10:@11215.4]
  assign _T_11162 = 4'h5 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11218.4]
  assign _T_11163 = _T_6208 & _T_11162; // @[LoadQueue.scala 131:72:@11219.4]
  assign _T_11165 = offsetQ_14 < 4'h5; // @[LoadQueue.scala 132:33:@11220.4]
  assign _T_11168 = _T_11165 & _T_6217; // @[LoadQueue.scala 132:41:@11222.4]
  assign _T_11170 = _T_11168 == 1'h0; // @[LoadQueue.scala 132:9:@11223.4]
  assign storesToCheck_14_5 = _T_2656 ? _T_11163 : _T_11170; // @[LoadQueue.scala 131:10:@11224.4]
  assign _T_11176 = 4'h6 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11227.4]
  assign _T_11177 = _T_6225 & _T_11176; // @[LoadQueue.scala 131:72:@11228.4]
  assign _T_11179 = offsetQ_14 < 4'h6; // @[LoadQueue.scala 132:33:@11229.4]
  assign _T_11182 = _T_11179 & _T_6234; // @[LoadQueue.scala 132:41:@11231.4]
  assign _T_11184 = _T_11182 == 1'h0; // @[LoadQueue.scala 132:9:@11232.4]
  assign storesToCheck_14_6 = _T_2656 ? _T_11177 : _T_11184; // @[LoadQueue.scala 131:10:@11233.4]
  assign _T_11190 = 4'h7 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11236.4]
  assign _T_11191 = _T_6242 & _T_11190; // @[LoadQueue.scala 131:72:@11237.4]
  assign _T_11193 = offsetQ_14 < 4'h7; // @[LoadQueue.scala 132:33:@11238.4]
  assign _T_11196 = _T_11193 & _T_6251; // @[LoadQueue.scala 132:41:@11240.4]
  assign _T_11198 = _T_11196 == 1'h0; // @[LoadQueue.scala 132:9:@11241.4]
  assign storesToCheck_14_7 = _T_2656 ? _T_11191 : _T_11198; // @[LoadQueue.scala 131:10:@11242.4]
  assign _T_11204 = 4'h8 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11245.4]
  assign _T_11205 = _T_6259 & _T_11204; // @[LoadQueue.scala 131:72:@11246.4]
  assign _T_11207 = offsetQ_14 < 4'h8; // @[LoadQueue.scala 132:33:@11247.4]
  assign _T_11210 = _T_11207 & _T_6268; // @[LoadQueue.scala 132:41:@11249.4]
  assign _T_11212 = _T_11210 == 1'h0; // @[LoadQueue.scala 132:9:@11250.4]
  assign storesToCheck_14_8 = _T_2656 ? _T_11205 : _T_11212; // @[LoadQueue.scala 131:10:@11251.4]
  assign _T_11218 = 4'h9 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11254.4]
  assign _T_11219 = _T_6276 & _T_11218; // @[LoadQueue.scala 131:72:@11255.4]
  assign _T_11221 = offsetQ_14 < 4'h9; // @[LoadQueue.scala 132:33:@11256.4]
  assign _T_11224 = _T_11221 & _T_6285; // @[LoadQueue.scala 132:41:@11258.4]
  assign _T_11226 = _T_11224 == 1'h0; // @[LoadQueue.scala 132:9:@11259.4]
  assign storesToCheck_14_9 = _T_2656 ? _T_11219 : _T_11226; // @[LoadQueue.scala 131:10:@11260.4]
  assign _T_11232 = 4'ha <= offsetQ_14; // @[LoadQueue.scala 131:81:@11263.4]
  assign _T_11233 = _T_6293 & _T_11232; // @[LoadQueue.scala 131:72:@11264.4]
  assign _T_11235 = offsetQ_14 < 4'ha; // @[LoadQueue.scala 132:33:@11265.4]
  assign _T_11238 = _T_11235 & _T_6302; // @[LoadQueue.scala 132:41:@11267.4]
  assign _T_11240 = _T_11238 == 1'h0; // @[LoadQueue.scala 132:9:@11268.4]
  assign storesToCheck_14_10 = _T_2656 ? _T_11233 : _T_11240; // @[LoadQueue.scala 131:10:@11269.4]
  assign _T_11246 = 4'hb <= offsetQ_14; // @[LoadQueue.scala 131:81:@11272.4]
  assign _T_11247 = _T_6310 & _T_11246; // @[LoadQueue.scala 131:72:@11273.4]
  assign _T_11249 = offsetQ_14 < 4'hb; // @[LoadQueue.scala 132:33:@11274.4]
  assign _T_11252 = _T_11249 & _T_6319; // @[LoadQueue.scala 132:41:@11276.4]
  assign _T_11254 = _T_11252 == 1'h0; // @[LoadQueue.scala 132:9:@11277.4]
  assign storesToCheck_14_11 = _T_2656 ? _T_11247 : _T_11254; // @[LoadQueue.scala 131:10:@11278.4]
  assign _T_11260 = 4'hc <= offsetQ_14; // @[LoadQueue.scala 131:81:@11281.4]
  assign _T_11261 = _T_6327 & _T_11260; // @[LoadQueue.scala 131:72:@11282.4]
  assign _T_11263 = offsetQ_14 < 4'hc; // @[LoadQueue.scala 132:33:@11283.4]
  assign _T_11266 = _T_11263 & _T_6336; // @[LoadQueue.scala 132:41:@11285.4]
  assign _T_11268 = _T_11266 == 1'h0; // @[LoadQueue.scala 132:9:@11286.4]
  assign storesToCheck_14_12 = _T_2656 ? _T_11261 : _T_11268; // @[LoadQueue.scala 131:10:@11287.4]
  assign _T_11274 = 4'hd <= offsetQ_14; // @[LoadQueue.scala 131:81:@11290.4]
  assign _T_11275 = _T_6344 & _T_11274; // @[LoadQueue.scala 131:72:@11291.4]
  assign _T_11277 = offsetQ_14 < 4'hd; // @[LoadQueue.scala 132:33:@11292.4]
  assign _T_11280 = _T_11277 & _T_6353; // @[LoadQueue.scala 132:41:@11294.4]
  assign _T_11282 = _T_11280 == 1'h0; // @[LoadQueue.scala 132:9:@11295.4]
  assign storesToCheck_14_13 = _T_2656 ? _T_11275 : _T_11282; // @[LoadQueue.scala 131:10:@11296.4]
  assign _T_11288 = 4'he <= offsetQ_14; // @[LoadQueue.scala 131:81:@11299.4]
  assign _T_11289 = _T_6361 & _T_11288; // @[LoadQueue.scala 131:72:@11300.4]
  assign _T_11291 = offsetQ_14 < 4'he; // @[LoadQueue.scala 132:33:@11301.4]
  assign _T_11294 = _T_11291 & _T_6370; // @[LoadQueue.scala 132:41:@11303.4]
  assign _T_11296 = _T_11294 == 1'h0; // @[LoadQueue.scala 132:9:@11304.4]
  assign storesToCheck_14_14 = _T_2656 ? _T_11289 : _T_11296; // @[LoadQueue.scala 131:10:@11305.4]
  assign _T_11302 = 4'hf <= offsetQ_14; // @[LoadQueue.scala 131:81:@11308.4]
  assign storesToCheck_14_15 = _T_2656 ? _T_11302 : 1'h1; // @[LoadQueue.scala 131:10:@11314.4]
  assign storesToCheck_15_0 = _T_2686 ? _T_6123 : 1'h1; // @[LoadQueue.scala 131:10:@11356.4]
  assign _T_11352 = 4'h1 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11359.4]
  assign _T_11353 = _T_6140 & _T_11352; // @[LoadQueue.scala 131:72:@11360.4]
  assign _T_11355 = offsetQ_15 < 4'h1; // @[LoadQueue.scala 132:33:@11361.4]
  assign _T_11358 = _T_11355 & _T_6149; // @[LoadQueue.scala 132:41:@11363.4]
  assign _T_11360 = _T_11358 == 1'h0; // @[LoadQueue.scala 132:9:@11364.4]
  assign storesToCheck_15_1 = _T_2686 ? _T_11353 : _T_11360; // @[LoadQueue.scala 131:10:@11365.4]
  assign _T_11366 = 4'h2 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11368.4]
  assign _T_11367 = _T_6157 & _T_11366; // @[LoadQueue.scala 131:72:@11369.4]
  assign _T_11369 = offsetQ_15 < 4'h2; // @[LoadQueue.scala 132:33:@11370.4]
  assign _T_11372 = _T_11369 & _T_6166; // @[LoadQueue.scala 132:41:@11372.4]
  assign _T_11374 = _T_11372 == 1'h0; // @[LoadQueue.scala 132:9:@11373.4]
  assign storesToCheck_15_2 = _T_2686 ? _T_11367 : _T_11374; // @[LoadQueue.scala 131:10:@11374.4]
  assign _T_11380 = 4'h3 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11377.4]
  assign _T_11381 = _T_6174 & _T_11380; // @[LoadQueue.scala 131:72:@11378.4]
  assign _T_11383 = offsetQ_15 < 4'h3; // @[LoadQueue.scala 132:33:@11379.4]
  assign _T_11386 = _T_11383 & _T_6183; // @[LoadQueue.scala 132:41:@11381.4]
  assign _T_11388 = _T_11386 == 1'h0; // @[LoadQueue.scala 132:9:@11382.4]
  assign storesToCheck_15_3 = _T_2686 ? _T_11381 : _T_11388; // @[LoadQueue.scala 131:10:@11383.4]
  assign _T_11394 = 4'h4 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11386.4]
  assign _T_11395 = _T_6191 & _T_11394; // @[LoadQueue.scala 131:72:@11387.4]
  assign _T_11397 = offsetQ_15 < 4'h4; // @[LoadQueue.scala 132:33:@11388.4]
  assign _T_11400 = _T_11397 & _T_6200; // @[LoadQueue.scala 132:41:@11390.4]
  assign _T_11402 = _T_11400 == 1'h0; // @[LoadQueue.scala 132:9:@11391.4]
  assign storesToCheck_15_4 = _T_2686 ? _T_11395 : _T_11402; // @[LoadQueue.scala 131:10:@11392.4]
  assign _T_11408 = 4'h5 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11395.4]
  assign _T_11409 = _T_6208 & _T_11408; // @[LoadQueue.scala 131:72:@11396.4]
  assign _T_11411 = offsetQ_15 < 4'h5; // @[LoadQueue.scala 132:33:@11397.4]
  assign _T_11414 = _T_11411 & _T_6217; // @[LoadQueue.scala 132:41:@11399.4]
  assign _T_11416 = _T_11414 == 1'h0; // @[LoadQueue.scala 132:9:@11400.4]
  assign storesToCheck_15_5 = _T_2686 ? _T_11409 : _T_11416; // @[LoadQueue.scala 131:10:@11401.4]
  assign _T_11422 = 4'h6 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11404.4]
  assign _T_11423 = _T_6225 & _T_11422; // @[LoadQueue.scala 131:72:@11405.4]
  assign _T_11425 = offsetQ_15 < 4'h6; // @[LoadQueue.scala 132:33:@11406.4]
  assign _T_11428 = _T_11425 & _T_6234; // @[LoadQueue.scala 132:41:@11408.4]
  assign _T_11430 = _T_11428 == 1'h0; // @[LoadQueue.scala 132:9:@11409.4]
  assign storesToCheck_15_6 = _T_2686 ? _T_11423 : _T_11430; // @[LoadQueue.scala 131:10:@11410.4]
  assign _T_11436 = 4'h7 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11413.4]
  assign _T_11437 = _T_6242 & _T_11436; // @[LoadQueue.scala 131:72:@11414.4]
  assign _T_11439 = offsetQ_15 < 4'h7; // @[LoadQueue.scala 132:33:@11415.4]
  assign _T_11442 = _T_11439 & _T_6251; // @[LoadQueue.scala 132:41:@11417.4]
  assign _T_11444 = _T_11442 == 1'h0; // @[LoadQueue.scala 132:9:@11418.4]
  assign storesToCheck_15_7 = _T_2686 ? _T_11437 : _T_11444; // @[LoadQueue.scala 131:10:@11419.4]
  assign _T_11450 = 4'h8 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11422.4]
  assign _T_11451 = _T_6259 & _T_11450; // @[LoadQueue.scala 131:72:@11423.4]
  assign _T_11453 = offsetQ_15 < 4'h8; // @[LoadQueue.scala 132:33:@11424.4]
  assign _T_11456 = _T_11453 & _T_6268; // @[LoadQueue.scala 132:41:@11426.4]
  assign _T_11458 = _T_11456 == 1'h0; // @[LoadQueue.scala 132:9:@11427.4]
  assign storesToCheck_15_8 = _T_2686 ? _T_11451 : _T_11458; // @[LoadQueue.scala 131:10:@11428.4]
  assign _T_11464 = 4'h9 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11431.4]
  assign _T_11465 = _T_6276 & _T_11464; // @[LoadQueue.scala 131:72:@11432.4]
  assign _T_11467 = offsetQ_15 < 4'h9; // @[LoadQueue.scala 132:33:@11433.4]
  assign _T_11470 = _T_11467 & _T_6285; // @[LoadQueue.scala 132:41:@11435.4]
  assign _T_11472 = _T_11470 == 1'h0; // @[LoadQueue.scala 132:9:@11436.4]
  assign storesToCheck_15_9 = _T_2686 ? _T_11465 : _T_11472; // @[LoadQueue.scala 131:10:@11437.4]
  assign _T_11478 = 4'ha <= offsetQ_15; // @[LoadQueue.scala 131:81:@11440.4]
  assign _T_11479 = _T_6293 & _T_11478; // @[LoadQueue.scala 131:72:@11441.4]
  assign _T_11481 = offsetQ_15 < 4'ha; // @[LoadQueue.scala 132:33:@11442.4]
  assign _T_11484 = _T_11481 & _T_6302; // @[LoadQueue.scala 132:41:@11444.4]
  assign _T_11486 = _T_11484 == 1'h0; // @[LoadQueue.scala 132:9:@11445.4]
  assign storesToCheck_15_10 = _T_2686 ? _T_11479 : _T_11486; // @[LoadQueue.scala 131:10:@11446.4]
  assign _T_11492 = 4'hb <= offsetQ_15; // @[LoadQueue.scala 131:81:@11449.4]
  assign _T_11493 = _T_6310 & _T_11492; // @[LoadQueue.scala 131:72:@11450.4]
  assign _T_11495 = offsetQ_15 < 4'hb; // @[LoadQueue.scala 132:33:@11451.4]
  assign _T_11498 = _T_11495 & _T_6319; // @[LoadQueue.scala 132:41:@11453.4]
  assign _T_11500 = _T_11498 == 1'h0; // @[LoadQueue.scala 132:9:@11454.4]
  assign storesToCheck_15_11 = _T_2686 ? _T_11493 : _T_11500; // @[LoadQueue.scala 131:10:@11455.4]
  assign _T_11506 = 4'hc <= offsetQ_15; // @[LoadQueue.scala 131:81:@11458.4]
  assign _T_11507 = _T_6327 & _T_11506; // @[LoadQueue.scala 131:72:@11459.4]
  assign _T_11509 = offsetQ_15 < 4'hc; // @[LoadQueue.scala 132:33:@11460.4]
  assign _T_11512 = _T_11509 & _T_6336; // @[LoadQueue.scala 132:41:@11462.4]
  assign _T_11514 = _T_11512 == 1'h0; // @[LoadQueue.scala 132:9:@11463.4]
  assign storesToCheck_15_12 = _T_2686 ? _T_11507 : _T_11514; // @[LoadQueue.scala 131:10:@11464.4]
  assign _T_11520 = 4'hd <= offsetQ_15; // @[LoadQueue.scala 131:81:@11467.4]
  assign _T_11521 = _T_6344 & _T_11520; // @[LoadQueue.scala 131:72:@11468.4]
  assign _T_11523 = offsetQ_15 < 4'hd; // @[LoadQueue.scala 132:33:@11469.4]
  assign _T_11526 = _T_11523 & _T_6353; // @[LoadQueue.scala 132:41:@11471.4]
  assign _T_11528 = _T_11526 == 1'h0; // @[LoadQueue.scala 132:9:@11472.4]
  assign storesToCheck_15_13 = _T_2686 ? _T_11521 : _T_11528; // @[LoadQueue.scala 131:10:@11473.4]
  assign _T_11534 = 4'he <= offsetQ_15; // @[LoadQueue.scala 131:81:@11476.4]
  assign _T_11535 = _T_6361 & _T_11534; // @[LoadQueue.scala 131:72:@11477.4]
  assign _T_11537 = offsetQ_15 < 4'he; // @[LoadQueue.scala 132:33:@11478.4]
  assign _T_11540 = _T_11537 & _T_6370; // @[LoadQueue.scala 132:41:@11480.4]
  assign _T_11542 = _T_11540 == 1'h0; // @[LoadQueue.scala 132:9:@11481.4]
  assign storesToCheck_15_14 = _T_2686 ? _T_11535 : _T_11542; // @[LoadQueue.scala 131:10:@11482.4]
  assign _T_11548 = 4'hf <= offsetQ_15; // @[LoadQueue.scala 131:81:@11485.4]
  assign storesToCheck_15_15 = _T_2686 ? _T_11548 : 1'h1; // @[LoadQueue.scala 131:10:@11491.4]
  assign _T_12810 = storesToCheck_0_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11526.4]
  assign entriesToCheck_0_0 = _T_12810 & checkBits_0; // @[LoadQueue.scala 141:26:@11527.4]
  assign _T_12812 = storesToCheck_0_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11528.4]
  assign entriesToCheck_0_1 = _T_12812 & checkBits_0; // @[LoadQueue.scala 141:26:@11529.4]
  assign _T_12814 = storesToCheck_0_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11530.4]
  assign entriesToCheck_0_2 = _T_12814 & checkBits_0; // @[LoadQueue.scala 141:26:@11531.4]
  assign _T_12816 = storesToCheck_0_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11532.4]
  assign entriesToCheck_0_3 = _T_12816 & checkBits_0; // @[LoadQueue.scala 141:26:@11533.4]
  assign _T_12818 = storesToCheck_0_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11534.4]
  assign entriesToCheck_0_4 = _T_12818 & checkBits_0; // @[LoadQueue.scala 141:26:@11535.4]
  assign _T_12820 = storesToCheck_0_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11536.4]
  assign entriesToCheck_0_5 = _T_12820 & checkBits_0; // @[LoadQueue.scala 141:26:@11537.4]
  assign _T_12822 = storesToCheck_0_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11538.4]
  assign entriesToCheck_0_6 = _T_12822 & checkBits_0; // @[LoadQueue.scala 141:26:@11539.4]
  assign _T_12824 = storesToCheck_0_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11540.4]
  assign entriesToCheck_0_7 = _T_12824 & checkBits_0; // @[LoadQueue.scala 141:26:@11541.4]
  assign _T_12826 = storesToCheck_0_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11542.4]
  assign entriesToCheck_0_8 = _T_12826 & checkBits_0; // @[LoadQueue.scala 141:26:@11543.4]
  assign _T_12828 = storesToCheck_0_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11544.4]
  assign entriesToCheck_0_9 = _T_12828 & checkBits_0; // @[LoadQueue.scala 141:26:@11545.4]
  assign _T_12830 = storesToCheck_0_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11546.4]
  assign entriesToCheck_0_10 = _T_12830 & checkBits_0; // @[LoadQueue.scala 141:26:@11547.4]
  assign _T_12832 = storesToCheck_0_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11548.4]
  assign entriesToCheck_0_11 = _T_12832 & checkBits_0; // @[LoadQueue.scala 141:26:@11549.4]
  assign _T_12834 = storesToCheck_0_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11550.4]
  assign entriesToCheck_0_12 = _T_12834 & checkBits_0; // @[LoadQueue.scala 141:26:@11551.4]
  assign _T_12836 = storesToCheck_0_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11552.4]
  assign entriesToCheck_0_13 = _T_12836 & checkBits_0; // @[LoadQueue.scala 141:26:@11553.4]
  assign _T_12838 = storesToCheck_0_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11554.4]
  assign entriesToCheck_0_14 = _T_12838 & checkBits_0; // @[LoadQueue.scala 141:26:@11555.4]
  assign _T_12840 = storesToCheck_0_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11556.4]
  assign entriesToCheck_0_15 = _T_12840 & checkBits_0; // @[LoadQueue.scala 141:26:@11557.4]
  assign _T_12842 = storesToCheck_1_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11574.4]
  assign entriesToCheck_1_0 = _T_12842 & checkBits_1; // @[LoadQueue.scala 141:26:@11575.4]
  assign _T_12844 = storesToCheck_1_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11576.4]
  assign entriesToCheck_1_1 = _T_12844 & checkBits_1; // @[LoadQueue.scala 141:26:@11577.4]
  assign _T_12846 = storesToCheck_1_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11578.4]
  assign entriesToCheck_1_2 = _T_12846 & checkBits_1; // @[LoadQueue.scala 141:26:@11579.4]
  assign _T_12848 = storesToCheck_1_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11580.4]
  assign entriesToCheck_1_3 = _T_12848 & checkBits_1; // @[LoadQueue.scala 141:26:@11581.4]
  assign _T_12850 = storesToCheck_1_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11582.4]
  assign entriesToCheck_1_4 = _T_12850 & checkBits_1; // @[LoadQueue.scala 141:26:@11583.4]
  assign _T_12852 = storesToCheck_1_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11584.4]
  assign entriesToCheck_1_5 = _T_12852 & checkBits_1; // @[LoadQueue.scala 141:26:@11585.4]
  assign _T_12854 = storesToCheck_1_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11586.4]
  assign entriesToCheck_1_6 = _T_12854 & checkBits_1; // @[LoadQueue.scala 141:26:@11587.4]
  assign _T_12856 = storesToCheck_1_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11588.4]
  assign entriesToCheck_1_7 = _T_12856 & checkBits_1; // @[LoadQueue.scala 141:26:@11589.4]
  assign _T_12858 = storesToCheck_1_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11590.4]
  assign entriesToCheck_1_8 = _T_12858 & checkBits_1; // @[LoadQueue.scala 141:26:@11591.4]
  assign _T_12860 = storesToCheck_1_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11592.4]
  assign entriesToCheck_1_9 = _T_12860 & checkBits_1; // @[LoadQueue.scala 141:26:@11593.4]
  assign _T_12862 = storesToCheck_1_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11594.4]
  assign entriesToCheck_1_10 = _T_12862 & checkBits_1; // @[LoadQueue.scala 141:26:@11595.4]
  assign _T_12864 = storesToCheck_1_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11596.4]
  assign entriesToCheck_1_11 = _T_12864 & checkBits_1; // @[LoadQueue.scala 141:26:@11597.4]
  assign _T_12866 = storesToCheck_1_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11598.4]
  assign entriesToCheck_1_12 = _T_12866 & checkBits_1; // @[LoadQueue.scala 141:26:@11599.4]
  assign _T_12868 = storesToCheck_1_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11600.4]
  assign entriesToCheck_1_13 = _T_12868 & checkBits_1; // @[LoadQueue.scala 141:26:@11601.4]
  assign _T_12870 = storesToCheck_1_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11602.4]
  assign entriesToCheck_1_14 = _T_12870 & checkBits_1; // @[LoadQueue.scala 141:26:@11603.4]
  assign _T_12872 = storesToCheck_1_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11604.4]
  assign entriesToCheck_1_15 = _T_12872 & checkBits_1; // @[LoadQueue.scala 141:26:@11605.4]
  assign _T_12874 = storesToCheck_2_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11622.4]
  assign entriesToCheck_2_0 = _T_12874 & checkBits_2; // @[LoadQueue.scala 141:26:@11623.4]
  assign _T_12876 = storesToCheck_2_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11624.4]
  assign entriesToCheck_2_1 = _T_12876 & checkBits_2; // @[LoadQueue.scala 141:26:@11625.4]
  assign _T_12878 = storesToCheck_2_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11626.4]
  assign entriesToCheck_2_2 = _T_12878 & checkBits_2; // @[LoadQueue.scala 141:26:@11627.4]
  assign _T_12880 = storesToCheck_2_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11628.4]
  assign entriesToCheck_2_3 = _T_12880 & checkBits_2; // @[LoadQueue.scala 141:26:@11629.4]
  assign _T_12882 = storesToCheck_2_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11630.4]
  assign entriesToCheck_2_4 = _T_12882 & checkBits_2; // @[LoadQueue.scala 141:26:@11631.4]
  assign _T_12884 = storesToCheck_2_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11632.4]
  assign entriesToCheck_2_5 = _T_12884 & checkBits_2; // @[LoadQueue.scala 141:26:@11633.4]
  assign _T_12886 = storesToCheck_2_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11634.4]
  assign entriesToCheck_2_6 = _T_12886 & checkBits_2; // @[LoadQueue.scala 141:26:@11635.4]
  assign _T_12888 = storesToCheck_2_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11636.4]
  assign entriesToCheck_2_7 = _T_12888 & checkBits_2; // @[LoadQueue.scala 141:26:@11637.4]
  assign _T_12890 = storesToCheck_2_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11638.4]
  assign entriesToCheck_2_8 = _T_12890 & checkBits_2; // @[LoadQueue.scala 141:26:@11639.4]
  assign _T_12892 = storesToCheck_2_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11640.4]
  assign entriesToCheck_2_9 = _T_12892 & checkBits_2; // @[LoadQueue.scala 141:26:@11641.4]
  assign _T_12894 = storesToCheck_2_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11642.4]
  assign entriesToCheck_2_10 = _T_12894 & checkBits_2; // @[LoadQueue.scala 141:26:@11643.4]
  assign _T_12896 = storesToCheck_2_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11644.4]
  assign entriesToCheck_2_11 = _T_12896 & checkBits_2; // @[LoadQueue.scala 141:26:@11645.4]
  assign _T_12898 = storesToCheck_2_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11646.4]
  assign entriesToCheck_2_12 = _T_12898 & checkBits_2; // @[LoadQueue.scala 141:26:@11647.4]
  assign _T_12900 = storesToCheck_2_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11648.4]
  assign entriesToCheck_2_13 = _T_12900 & checkBits_2; // @[LoadQueue.scala 141:26:@11649.4]
  assign _T_12902 = storesToCheck_2_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11650.4]
  assign entriesToCheck_2_14 = _T_12902 & checkBits_2; // @[LoadQueue.scala 141:26:@11651.4]
  assign _T_12904 = storesToCheck_2_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11652.4]
  assign entriesToCheck_2_15 = _T_12904 & checkBits_2; // @[LoadQueue.scala 141:26:@11653.4]
  assign _T_12906 = storesToCheck_3_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11670.4]
  assign entriesToCheck_3_0 = _T_12906 & checkBits_3; // @[LoadQueue.scala 141:26:@11671.4]
  assign _T_12908 = storesToCheck_3_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11672.4]
  assign entriesToCheck_3_1 = _T_12908 & checkBits_3; // @[LoadQueue.scala 141:26:@11673.4]
  assign _T_12910 = storesToCheck_3_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11674.4]
  assign entriesToCheck_3_2 = _T_12910 & checkBits_3; // @[LoadQueue.scala 141:26:@11675.4]
  assign _T_12912 = storesToCheck_3_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11676.4]
  assign entriesToCheck_3_3 = _T_12912 & checkBits_3; // @[LoadQueue.scala 141:26:@11677.4]
  assign _T_12914 = storesToCheck_3_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11678.4]
  assign entriesToCheck_3_4 = _T_12914 & checkBits_3; // @[LoadQueue.scala 141:26:@11679.4]
  assign _T_12916 = storesToCheck_3_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11680.4]
  assign entriesToCheck_3_5 = _T_12916 & checkBits_3; // @[LoadQueue.scala 141:26:@11681.4]
  assign _T_12918 = storesToCheck_3_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11682.4]
  assign entriesToCheck_3_6 = _T_12918 & checkBits_3; // @[LoadQueue.scala 141:26:@11683.4]
  assign _T_12920 = storesToCheck_3_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11684.4]
  assign entriesToCheck_3_7 = _T_12920 & checkBits_3; // @[LoadQueue.scala 141:26:@11685.4]
  assign _T_12922 = storesToCheck_3_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11686.4]
  assign entriesToCheck_3_8 = _T_12922 & checkBits_3; // @[LoadQueue.scala 141:26:@11687.4]
  assign _T_12924 = storesToCheck_3_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11688.4]
  assign entriesToCheck_3_9 = _T_12924 & checkBits_3; // @[LoadQueue.scala 141:26:@11689.4]
  assign _T_12926 = storesToCheck_3_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11690.4]
  assign entriesToCheck_3_10 = _T_12926 & checkBits_3; // @[LoadQueue.scala 141:26:@11691.4]
  assign _T_12928 = storesToCheck_3_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11692.4]
  assign entriesToCheck_3_11 = _T_12928 & checkBits_3; // @[LoadQueue.scala 141:26:@11693.4]
  assign _T_12930 = storesToCheck_3_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11694.4]
  assign entriesToCheck_3_12 = _T_12930 & checkBits_3; // @[LoadQueue.scala 141:26:@11695.4]
  assign _T_12932 = storesToCheck_3_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11696.4]
  assign entriesToCheck_3_13 = _T_12932 & checkBits_3; // @[LoadQueue.scala 141:26:@11697.4]
  assign _T_12934 = storesToCheck_3_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11698.4]
  assign entriesToCheck_3_14 = _T_12934 & checkBits_3; // @[LoadQueue.scala 141:26:@11699.4]
  assign _T_12936 = storesToCheck_3_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11700.4]
  assign entriesToCheck_3_15 = _T_12936 & checkBits_3; // @[LoadQueue.scala 141:26:@11701.4]
  assign _T_12938 = storesToCheck_4_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11718.4]
  assign entriesToCheck_4_0 = _T_12938 & checkBits_4; // @[LoadQueue.scala 141:26:@11719.4]
  assign _T_12940 = storesToCheck_4_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11720.4]
  assign entriesToCheck_4_1 = _T_12940 & checkBits_4; // @[LoadQueue.scala 141:26:@11721.4]
  assign _T_12942 = storesToCheck_4_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11722.4]
  assign entriesToCheck_4_2 = _T_12942 & checkBits_4; // @[LoadQueue.scala 141:26:@11723.4]
  assign _T_12944 = storesToCheck_4_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11724.4]
  assign entriesToCheck_4_3 = _T_12944 & checkBits_4; // @[LoadQueue.scala 141:26:@11725.4]
  assign _T_12946 = storesToCheck_4_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11726.4]
  assign entriesToCheck_4_4 = _T_12946 & checkBits_4; // @[LoadQueue.scala 141:26:@11727.4]
  assign _T_12948 = storesToCheck_4_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11728.4]
  assign entriesToCheck_4_5 = _T_12948 & checkBits_4; // @[LoadQueue.scala 141:26:@11729.4]
  assign _T_12950 = storesToCheck_4_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11730.4]
  assign entriesToCheck_4_6 = _T_12950 & checkBits_4; // @[LoadQueue.scala 141:26:@11731.4]
  assign _T_12952 = storesToCheck_4_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11732.4]
  assign entriesToCheck_4_7 = _T_12952 & checkBits_4; // @[LoadQueue.scala 141:26:@11733.4]
  assign _T_12954 = storesToCheck_4_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11734.4]
  assign entriesToCheck_4_8 = _T_12954 & checkBits_4; // @[LoadQueue.scala 141:26:@11735.4]
  assign _T_12956 = storesToCheck_4_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11736.4]
  assign entriesToCheck_4_9 = _T_12956 & checkBits_4; // @[LoadQueue.scala 141:26:@11737.4]
  assign _T_12958 = storesToCheck_4_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11738.4]
  assign entriesToCheck_4_10 = _T_12958 & checkBits_4; // @[LoadQueue.scala 141:26:@11739.4]
  assign _T_12960 = storesToCheck_4_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11740.4]
  assign entriesToCheck_4_11 = _T_12960 & checkBits_4; // @[LoadQueue.scala 141:26:@11741.4]
  assign _T_12962 = storesToCheck_4_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11742.4]
  assign entriesToCheck_4_12 = _T_12962 & checkBits_4; // @[LoadQueue.scala 141:26:@11743.4]
  assign _T_12964 = storesToCheck_4_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11744.4]
  assign entriesToCheck_4_13 = _T_12964 & checkBits_4; // @[LoadQueue.scala 141:26:@11745.4]
  assign _T_12966 = storesToCheck_4_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11746.4]
  assign entriesToCheck_4_14 = _T_12966 & checkBits_4; // @[LoadQueue.scala 141:26:@11747.4]
  assign _T_12968 = storesToCheck_4_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11748.4]
  assign entriesToCheck_4_15 = _T_12968 & checkBits_4; // @[LoadQueue.scala 141:26:@11749.4]
  assign _T_12970 = storesToCheck_5_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11766.4]
  assign entriesToCheck_5_0 = _T_12970 & checkBits_5; // @[LoadQueue.scala 141:26:@11767.4]
  assign _T_12972 = storesToCheck_5_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11768.4]
  assign entriesToCheck_5_1 = _T_12972 & checkBits_5; // @[LoadQueue.scala 141:26:@11769.4]
  assign _T_12974 = storesToCheck_5_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11770.4]
  assign entriesToCheck_5_2 = _T_12974 & checkBits_5; // @[LoadQueue.scala 141:26:@11771.4]
  assign _T_12976 = storesToCheck_5_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11772.4]
  assign entriesToCheck_5_3 = _T_12976 & checkBits_5; // @[LoadQueue.scala 141:26:@11773.4]
  assign _T_12978 = storesToCheck_5_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11774.4]
  assign entriesToCheck_5_4 = _T_12978 & checkBits_5; // @[LoadQueue.scala 141:26:@11775.4]
  assign _T_12980 = storesToCheck_5_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11776.4]
  assign entriesToCheck_5_5 = _T_12980 & checkBits_5; // @[LoadQueue.scala 141:26:@11777.4]
  assign _T_12982 = storesToCheck_5_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11778.4]
  assign entriesToCheck_5_6 = _T_12982 & checkBits_5; // @[LoadQueue.scala 141:26:@11779.4]
  assign _T_12984 = storesToCheck_5_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11780.4]
  assign entriesToCheck_5_7 = _T_12984 & checkBits_5; // @[LoadQueue.scala 141:26:@11781.4]
  assign _T_12986 = storesToCheck_5_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11782.4]
  assign entriesToCheck_5_8 = _T_12986 & checkBits_5; // @[LoadQueue.scala 141:26:@11783.4]
  assign _T_12988 = storesToCheck_5_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11784.4]
  assign entriesToCheck_5_9 = _T_12988 & checkBits_5; // @[LoadQueue.scala 141:26:@11785.4]
  assign _T_12990 = storesToCheck_5_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11786.4]
  assign entriesToCheck_5_10 = _T_12990 & checkBits_5; // @[LoadQueue.scala 141:26:@11787.4]
  assign _T_12992 = storesToCheck_5_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11788.4]
  assign entriesToCheck_5_11 = _T_12992 & checkBits_5; // @[LoadQueue.scala 141:26:@11789.4]
  assign _T_12994 = storesToCheck_5_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11790.4]
  assign entriesToCheck_5_12 = _T_12994 & checkBits_5; // @[LoadQueue.scala 141:26:@11791.4]
  assign _T_12996 = storesToCheck_5_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11792.4]
  assign entriesToCheck_5_13 = _T_12996 & checkBits_5; // @[LoadQueue.scala 141:26:@11793.4]
  assign _T_12998 = storesToCheck_5_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11794.4]
  assign entriesToCheck_5_14 = _T_12998 & checkBits_5; // @[LoadQueue.scala 141:26:@11795.4]
  assign _T_13000 = storesToCheck_5_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11796.4]
  assign entriesToCheck_5_15 = _T_13000 & checkBits_5; // @[LoadQueue.scala 141:26:@11797.4]
  assign _T_13002 = storesToCheck_6_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11814.4]
  assign entriesToCheck_6_0 = _T_13002 & checkBits_6; // @[LoadQueue.scala 141:26:@11815.4]
  assign _T_13004 = storesToCheck_6_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11816.4]
  assign entriesToCheck_6_1 = _T_13004 & checkBits_6; // @[LoadQueue.scala 141:26:@11817.4]
  assign _T_13006 = storesToCheck_6_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11818.4]
  assign entriesToCheck_6_2 = _T_13006 & checkBits_6; // @[LoadQueue.scala 141:26:@11819.4]
  assign _T_13008 = storesToCheck_6_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11820.4]
  assign entriesToCheck_6_3 = _T_13008 & checkBits_6; // @[LoadQueue.scala 141:26:@11821.4]
  assign _T_13010 = storesToCheck_6_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11822.4]
  assign entriesToCheck_6_4 = _T_13010 & checkBits_6; // @[LoadQueue.scala 141:26:@11823.4]
  assign _T_13012 = storesToCheck_6_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11824.4]
  assign entriesToCheck_6_5 = _T_13012 & checkBits_6; // @[LoadQueue.scala 141:26:@11825.4]
  assign _T_13014 = storesToCheck_6_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11826.4]
  assign entriesToCheck_6_6 = _T_13014 & checkBits_6; // @[LoadQueue.scala 141:26:@11827.4]
  assign _T_13016 = storesToCheck_6_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11828.4]
  assign entriesToCheck_6_7 = _T_13016 & checkBits_6; // @[LoadQueue.scala 141:26:@11829.4]
  assign _T_13018 = storesToCheck_6_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11830.4]
  assign entriesToCheck_6_8 = _T_13018 & checkBits_6; // @[LoadQueue.scala 141:26:@11831.4]
  assign _T_13020 = storesToCheck_6_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11832.4]
  assign entriesToCheck_6_9 = _T_13020 & checkBits_6; // @[LoadQueue.scala 141:26:@11833.4]
  assign _T_13022 = storesToCheck_6_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11834.4]
  assign entriesToCheck_6_10 = _T_13022 & checkBits_6; // @[LoadQueue.scala 141:26:@11835.4]
  assign _T_13024 = storesToCheck_6_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11836.4]
  assign entriesToCheck_6_11 = _T_13024 & checkBits_6; // @[LoadQueue.scala 141:26:@11837.4]
  assign _T_13026 = storesToCheck_6_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11838.4]
  assign entriesToCheck_6_12 = _T_13026 & checkBits_6; // @[LoadQueue.scala 141:26:@11839.4]
  assign _T_13028 = storesToCheck_6_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11840.4]
  assign entriesToCheck_6_13 = _T_13028 & checkBits_6; // @[LoadQueue.scala 141:26:@11841.4]
  assign _T_13030 = storesToCheck_6_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11842.4]
  assign entriesToCheck_6_14 = _T_13030 & checkBits_6; // @[LoadQueue.scala 141:26:@11843.4]
  assign _T_13032 = storesToCheck_6_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11844.4]
  assign entriesToCheck_6_15 = _T_13032 & checkBits_6; // @[LoadQueue.scala 141:26:@11845.4]
  assign _T_13034 = storesToCheck_7_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11862.4]
  assign entriesToCheck_7_0 = _T_13034 & checkBits_7; // @[LoadQueue.scala 141:26:@11863.4]
  assign _T_13036 = storesToCheck_7_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11864.4]
  assign entriesToCheck_7_1 = _T_13036 & checkBits_7; // @[LoadQueue.scala 141:26:@11865.4]
  assign _T_13038 = storesToCheck_7_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11866.4]
  assign entriesToCheck_7_2 = _T_13038 & checkBits_7; // @[LoadQueue.scala 141:26:@11867.4]
  assign _T_13040 = storesToCheck_7_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11868.4]
  assign entriesToCheck_7_3 = _T_13040 & checkBits_7; // @[LoadQueue.scala 141:26:@11869.4]
  assign _T_13042 = storesToCheck_7_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11870.4]
  assign entriesToCheck_7_4 = _T_13042 & checkBits_7; // @[LoadQueue.scala 141:26:@11871.4]
  assign _T_13044 = storesToCheck_7_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11872.4]
  assign entriesToCheck_7_5 = _T_13044 & checkBits_7; // @[LoadQueue.scala 141:26:@11873.4]
  assign _T_13046 = storesToCheck_7_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11874.4]
  assign entriesToCheck_7_6 = _T_13046 & checkBits_7; // @[LoadQueue.scala 141:26:@11875.4]
  assign _T_13048 = storesToCheck_7_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11876.4]
  assign entriesToCheck_7_7 = _T_13048 & checkBits_7; // @[LoadQueue.scala 141:26:@11877.4]
  assign _T_13050 = storesToCheck_7_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11878.4]
  assign entriesToCheck_7_8 = _T_13050 & checkBits_7; // @[LoadQueue.scala 141:26:@11879.4]
  assign _T_13052 = storesToCheck_7_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11880.4]
  assign entriesToCheck_7_9 = _T_13052 & checkBits_7; // @[LoadQueue.scala 141:26:@11881.4]
  assign _T_13054 = storesToCheck_7_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11882.4]
  assign entriesToCheck_7_10 = _T_13054 & checkBits_7; // @[LoadQueue.scala 141:26:@11883.4]
  assign _T_13056 = storesToCheck_7_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11884.4]
  assign entriesToCheck_7_11 = _T_13056 & checkBits_7; // @[LoadQueue.scala 141:26:@11885.4]
  assign _T_13058 = storesToCheck_7_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11886.4]
  assign entriesToCheck_7_12 = _T_13058 & checkBits_7; // @[LoadQueue.scala 141:26:@11887.4]
  assign _T_13060 = storesToCheck_7_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11888.4]
  assign entriesToCheck_7_13 = _T_13060 & checkBits_7; // @[LoadQueue.scala 141:26:@11889.4]
  assign _T_13062 = storesToCheck_7_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11890.4]
  assign entriesToCheck_7_14 = _T_13062 & checkBits_7; // @[LoadQueue.scala 141:26:@11891.4]
  assign _T_13064 = storesToCheck_7_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11892.4]
  assign entriesToCheck_7_15 = _T_13064 & checkBits_7; // @[LoadQueue.scala 141:26:@11893.4]
  assign _T_13066 = storesToCheck_8_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11910.4]
  assign entriesToCheck_8_0 = _T_13066 & checkBits_8; // @[LoadQueue.scala 141:26:@11911.4]
  assign _T_13068 = storesToCheck_8_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11912.4]
  assign entriesToCheck_8_1 = _T_13068 & checkBits_8; // @[LoadQueue.scala 141:26:@11913.4]
  assign _T_13070 = storesToCheck_8_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11914.4]
  assign entriesToCheck_8_2 = _T_13070 & checkBits_8; // @[LoadQueue.scala 141:26:@11915.4]
  assign _T_13072 = storesToCheck_8_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11916.4]
  assign entriesToCheck_8_3 = _T_13072 & checkBits_8; // @[LoadQueue.scala 141:26:@11917.4]
  assign _T_13074 = storesToCheck_8_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11918.4]
  assign entriesToCheck_8_4 = _T_13074 & checkBits_8; // @[LoadQueue.scala 141:26:@11919.4]
  assign _T_13076 = storesToCheck_8_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11920.4]
  assign entriesToCheck_8_5 = _T_13076 & checkBits_8; // @[LoadQueue.scala 141:26:@11921.4]
  assign _T_13078 = storesToCheck_8_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11922.4]
  assign entriesToCheck_8_6 = _T_13078 & checkBits_8; // @[LoadQueue.scala 141:26:@11923.4]
  assign _T_13080 = storesToCheck_8_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11924.4]
  assign entriesToCheck_8_7 = _T_13080 & checkBits_8; // @[LoadQueue.scala 141:26:@11925.4]
  assign _T_13082 = storesToCheck_8_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11926.4]
  assign entriesToCheck_8_8 = _T_13082 & checkBits_8; // @[LoadQueue.scala 141:26:@11927.4]
  assign _T_13084 = storesToCheck_8_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11928.4]
  assign entriesToCheck_8_9 = _T_13084 & checkBits_8; // @[LoadQueue.scala 141:26:@11929.4]
  assign _T_13086 = storesToCheck_8_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11930.4]
  assign entriesToCheck_8_10 = _T_13086 & checkBits_8; // @[LoadQueue.scala 141:26:@11931.4]
  assign _T_13088 = storesToCheck_8_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11932.4]
  assign entriesToCheck_8_11 = _T_13088 & checkBits_8; // @[LoadQueue.scala 141:26:@11933.4]
  assign _T_13090 = storesToCheck_8_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11934.4]
  assign entriesToCheck_8_12 = _T_13090 & checkBits_8; // @[LoadQueue.scala 141:26:@11935.4]
  assign _T_13092 = storesToCheck_8_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11936.4]
  assign entriesToCheck_8_13 = _T_13092 & checkBits_8; // @[LoadQueue.scala 141:26:@11937.4]
  assign _T_13094 = storesToCheck_8_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11938.4]
  assign entriesToCheck_8_14 = _T_13094 & checkBits_8; // @[LoadQueue.scala 141:26:@11939.4]
  assign _T_13096 = storesToCheck_8_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11940.4]
  assign entriesToCheck_8_15 = _T_13096 & checkBits_8; // @[LoadQueue.scala 141:26:@11941.4]
  assign _T_13098 = storesToCheck_9_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11958.4]
  assign entriesToCheck_9_0 = _T_13098 & checkBits_9; // @[LoadQueue.scala 141:26:@11959.4]
  assign _T_13100 = storesToCheck_9_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11960.4]
  assign entriesToCheck_9_1 = _T_13100 & checkBits_9; // @[LoadQueue.scala 141:26:@11961.4]
  assign _T_13102 = storesToCheck_9_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11962.4]
  assign entriesToCheck_9_2 = _T_13102 & checkBits_9; // @[LoadQueue.scala 141:26:@11963.4]
  assign _T_13104 = storesToCheck_9_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11964.4]
  assign entriesToCheck_9_3 = _T_13104 & checkBits_9; // @[LoadQueue.scala 141:26:@11965.4]
  assign _T_13106 = storesToCheck_9_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11966.4]
  assign entriesToCheck_9_4 = _T_13106 & checkBits_9; // @[LoadQueue.scala 141:26:@11967.4]
  assign _T_13108 = storesToCheck_9_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11968.4]
  assign entriesToCheck_9_5 = _T_13108 & checkBits_9; // @[LoadQueue.scala 141:26:@11969.4]
  assign _T_13110 = storesToCheck_9_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11970.4]
  assign entriesToCheck_9_6 = _T_13110 & checkBits_9; // @[LoadQueue.scala 141:26:@11971.4]
  assign _T_13112 = storesToCheck_9_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11972.4]
  assign entriesToCheck_9_7 = _T_13112 & checkBits_9; // @[LoadQueue.scala 141:26:@11973.4]
  assign _T_13114 = storesToCheck_9_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11974.4]
  assign entriesToCheck_9_8 = _T_13114 & checkBits_9; // @[LoadQueue.scala 141:26:@11975.4]
  assign _T_13116 = storesToCheck_9_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11976.4]
  assign entriesToCheck_9_9 = _T_13116 & checkBits_9; // @[LoadQueue.scala 141:26:@11977.4]
  assign _T_13118 = storesToCheck_9_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11978.4]
  assign entriesToCheck_9_10 = _T_13118 & checkBits_9; // @[LoadQueue.scala 141:26:@11979.4]
  assign _T_13120 = storesToCheck_9_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11980.4]
  assign entriesToCheck_9_11 = _T_13120 & checkBits_9; // @[LoadQueue.scala 141:26:@11981.4]
  assign _T_13122 = storesToCheck_9_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11982.4]
  assign entriesToCheck_9_12 = _T_13122 & checkBits_9; // @[LoadQueue.scala 141:26:@11983.4]
  assign _T_13124 = storesToCheck_9_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11984.4]
  assign entriesToCheck_9_13 = _T_13124 & checkBits_9; // @[LoadQueue.scala 141:26:@11985.4]
  assign _T_13126 = storesToCheck_9_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11986.4]
  assign entriesToCheck_9_14 = _T_13126 & checkBits_9; // @[LoadQueue.scala 141:26:@11987.4]
  assign _T_13128 = storesToCheck_9_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11988.4]
  assign entriesToCheck_9_15 = _T_13128 & checkBits_9; // @[LoadQueue.scala 141:26:@11989.4]
  assign _T_13130 = storesToCheck_10_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@12006.4]
  assign entriesToCheck_10_0 = _T_13130 & checkBits_10; // @[LoadQueue.scala 141:26:@12007.4]
  assign _T_13132 = storesToCheck_10_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@12008.4]
  assign entriesToCheck_10_1 = _T_13132 & checkBits_10; // @[LoadQueue.scala 141:26:@12009.4]
  assign _T_13134 = storesToCheck_10_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@12010.4]
  assign entriesToCheck_10_2 = _T_13134 & checkBits_10; // @[LoadQueue.scala 141:26:@12011.4]
  assign _T_13136 = storesToCheck_10_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@12012.4]
  assign entriesToCheck_10_3 = _T_13136 & checkBits_10; // @[LoadQueue.scala 141:26:@12013.4]
  assign _T_13138 = storesToCheck_10_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@12014.4]
  assign entriesToCheck_10_4 = _T_13138 & checkBits_10; // @[LoadQueue.scala 141:26:@12015.4]
  assign _T_13140 = storesToCheck_10_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@12016.4]
  assign entriesToCheck_10_5 = _T_13140 & checkBits_10; // @[LoadQueue.scala 141:26:@12017.4]
  assign _T_13142 = storesToCheck_10_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@12018.4]
  assign entriesToCheck_10_6 = _T_13142 & checkBits_10; // @[LoadQueue.scala 141:26:@12019.4]
  assign _T_13144 = storesToCheck_10_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@12020.4]
  assign entriesToCheck_10_7 = _T_13144 & checkBits_10; // @[LoadQueue.scala 141:26:@12021.4]
  assign _T_13146 = storesToCheck_10_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@12022.4]
  assign entriesToCheck_10_8 = _T_13146 & checkBits_10; // @[LoadQueue.scala 141:26:@12023.4]
  assign _T_13148 = storesToCheck_10_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@12024.4]
  assign entriesToCheck_10_9 = _T_13148 & checkBits_10; // @[LoadQueue.scala 141:26:@12025.4]
  assign _T_13150 = storesToCheck_10_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@12026.4]
  assign entriesToCheck_10_10 = _T_13150 & checkBits_10; // @[LoadQueue.scala 141:26:@12027.4]
  assign _T_13152 = storesToCheck_10_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@12028.4]
  assign entriesToCheck_10_11 = _T_13152 & checkBits_10; // @[LoadQueue.scala 141:26:@12029.4]
  assign _T_13154 = storesToCheck_10_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@12030.4]
  assign entriesToCheck_10_12 = _T_13154 & checkBits_10; // @[LoadQueue.scala 141:26:@12031.4]
  assign _T_13156 = storesToCheck_10_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@12032.4]
  assign entriesToCheck_10_13 = _T_13156 & checkBits_10; // @[LoadQueue.scala 141:26:@12033.4]
  assign _T_13158 = storesToCheck_10_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@12034.4]
  assign entriesToCheck_10_14 = _T_13158 & checkBits_10; // @[LoadQueue.scala 141:26:@12035.4]
  assign _T_13160 = storesToCheck_10_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@12036.4]
  assign entriesToCheck_10_15 = _T_13160 & checkBits_10; // @[LoadQueue.scala 141:26:@12037.4]
  assign _T_13162 = storesToCheck_11_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@12054.4]
  assign entriesToCheck_11_0 = _T_13162 & checkBits_11; // @[LoadQueue.scala 141:26:@12055.4]
  assign _T_13164 = storesToCheck_11_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@12056.4]
  assign entriesToCheck_11_1 = _T_13164 & checkBits_11; // @[LoadQueue.scala 141:26:@12057.4]
  assign _T_13166 = storesToCheck_11_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@12058.4]
  assign entriesToCheck_11_2 = _T_13166 & checkBits_11; // @[LoadQueue.scala 141:26:@12059.4]
  assign _T_13168 = storesToCheck_11_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@12060.4]
  assign entriesToCheck_11_3 = _T_13168 & checkBits_11; // @[LoadQueue.scala 141:26:@12061.4]
  assign _T_13170 = storesToCheck_11_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@12062.4]
  assign entriesToCheck_11_4 = _T_13170 & checkBits_11; // @[LoadQueue.scala 141:26:@12063.4]
  assign _T_13172 = storesToCheck_11_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@12064.4]
  assign entriesToCheck_11_5 = _T_13172 & checkBits_11; // @[LoadQueue.scala 141:26:@12065.4]
  assign _T_13174 = storesToCheck_11_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@12066.4]
  assign entriesToCheck_11_6 = _T_13174 & checkBits_11; // @[LoadQueue.scala 141:26:@12067.4]
  assign _T_13176 = storesToCheck_11_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@12068.4]
  assign entriesToCheck_11_7 = _T_13176 & checkBits_11; // @[LoadQueue.scala 141:26:@12069.4]
  assign _T_13178 = storesToCheck_11_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@12070.4]
  assign entriesToCheck_11_8 = _T_13178 & checkBits_11; // @[LoadQueue.scala 141:26:@12071.4]
  assign _T_13180 = storesToCheck_11_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@12072.4]
  assign entriesToCheck_11_9 = _T_13180 & checkBits_11; // @[LoadQueue.scala 141:26:@12073.4]
  assign _T_13182 = storesToCheck_11_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@12074.4]
  assign entriesToCheck_11_10 = _T_13182 & checkBits_11; // @[LoadQueue.scala 141:26:@12075.4]
  assign _T_13184 = storesToCheck_11_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@12076.4]
  assign entriesToCheck_11_11 = _T_13184 & checkBits_11; // @[LoadQueue.scala 141:26:@12077.4]
  assign _T_13186 = storesToCheck_11_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@12078.4]
  assign entriesToCheck_11_12 = _T_13186 & checkBits_11; // @[LoadQueue.scala 141:26:@12079.4]
  assign _T_13188 = storesToCheck_11_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@12080.4]
  assign entriesToCheck_11_13 = _T_13188 & checkBits_11; // @[LoadQueue.scala 141:26:@12081.4]
  assign _T_13190 = storesToCheck_11_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@12082.4]
  assign entriesToCheck_11_14 = _T_13190 & checkBits_11; // @[LoadQueue.scala 141:26:@12083.4]
  assign _T_13192 = storesToCheck_11_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@12084.4]
  assign entriesToCheck_11_15 = _T_13192 & checkBits_11; // @[LoadQueue.scala 141:26:@12085.4]
  assign _T_13194 = storesToCheck_12_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@12102.4]
  assign entriesToCheck_12_0 = _T_13194 & checkBits_12; // @[LoadQueue.scala 141:26:@12103.4]
  assign _T_13196 = storesToCheck_12_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@12104.4]
  assign entriesToCheck_12_1 = _T_13196 & checkBits_12; // @[LoadQueue.scala 141:26:@12105.4]
  assign _T_13198 = storesToCheck_12_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@12106.4]
  assign entriesToCheck_12_2 = _T_13198 & checkBits_12; // @[LoadQueue.scala 141:26:@12107.4]
  assign _T_13200 = storesToCheck_12_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@12108.4]
  assign entriesToCheck_12_3 = _T_13200 & checkBits_12; // @[LoadQueue.scala 141:26:@12109.4]
  assign _T_13202 = storesToCheck_12_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@12110.4]
  assign entriesToCheck_12_4 = _T_13202 & checkBits_12; // @[LoadQueue.scala 141:26:@12111.4]
  assign _T_13204 = storesToCheck_12_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@12112.4]
  assign entriesToCheck_12_5 = _T_13204 & checkBits_12; // @[LoadQueue.scala 141:26:@12113.4]
  assign _T_13206 = storesToCheck_12_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@12114.4]
  assign entriesToCheck_12_6 = _T_13206 & checkBits_12; // @[LoadQueue.scala 141:26:@12115.4]
  assign _T_13208 = storesToCheck_12_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@12116.4]
  assign entriesToCheck_12_7 = _T_13208 & checkBits_12; // @[LoadQueue.scala 141:26:@12117.4]
  assign _T_13210 = storesToCheck_12_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@12118.4]
  assign entriesToCheck_12_8 = _T_13210 & checkBits_12; // @[LoadQueue.scala 141:26:@12119.4]
  assign _T_13212 = storesToCheck_12_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@12120.4]
  assign entriesToCheck_12_9 = _T_13212 & checkBits_12; // @[LoadQueue.scala 141:26:@12121.4]
  assign _T_13214 = storesToCheck_12_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@12122.4]
  assign entriesToCheck_12_10 = _T_13214 & checkBits_12; // @[LoadQueue.scala 141:26:@12123.4]
  assign _T_13216 = storesToCheck_12_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@12124.4]
  assign entriesToCheck_12_11 = _T_13216 & checkBits_12; // @[LoadQueue.scala 141:26:@12125.4]
  assign _T_13218 = storesToCheck_12_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@12126.4]
  assign entriesToCheck_12_12 = _T_13218 & checkBits_12; // @[LoadQueue.scala 141:26:@12127.4]
  assign _T_13220 = storesToCheck_12_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@12128.4]
  assign entriesToCheck_12_13 = _T_13220 & checkBits_12; // @[LoadQueue.scala 141:26:@12129.4]
  assign _T_13222 = storesToCheck_12_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@12130.4]
  assign entriesToCheck_12_14 = _T_13222 & checkBits_12; // @[LoadQueue.scala 141:26:@12131.4]
  assign _T_13224 = storesToCheck_12_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@12132.4]
  assign entriesToCheck_12_15 = _T_13224 & checkBits_12; // @[LoadQueue.scala 141:26:@12133.4]
  assign _T_13226 = storesToCheck_13_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@12150.4]
  assign entriesToCheck_13_0 = _T_13226 & checkBits_13; // @[LoadQueue.scala 141:26:@12151.4]
  assign _T_13228 = storesToCheck_13_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@12152.4]
  assign entriesToCheck_13_1 = _T_13228 & checkBits_13; // @[LoadQueue.scala 141:26:@12153.4]
  assign _T_13230 = storesToCheck_13_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@12154.4]
  assign entriesToCheck_13_2 = _T_13230 & checkBits_13; // @[LoadQueue.scala 141:26:@12155.4]
  assign _T_13232 = storesToCheck_13_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@12156.4]
  assign entriesToCheck_13_3 = _T_13232 & checkBits_13; // @[LoadQueue.scala 141:26:@12157.4]
  assign _T_13234 = storesToCheck_13_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@12158.4]
  assign entriesToCheck_13_4 = _T_13234 & checkBits_13; // @[LoadQueue.scala 141:26:@12159.4]
  assign _T_13236 = storesToCheck_13_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@12160.4]
  assign entriesToCheck_13_5 = _T_13236 & checkBits_13; // @[LoadQueue.scala 141:26:@12161.4]
  assign _T_13238 = storesToCheck_13_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@12162.4]
  assign entriesToCheck_13_6 = _T_13238 & checkBits_13; // @[LoadQueue.scala 141:26:@12163.4]
  assign _T_13240 = storesToCheck_13_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@12164.4]
  assign entriesToCheck_13_7 = _T_13240 & checkBits_13; // @[LoadQueue.scala 141:26:@12165.4]
  assign _T_13242 = storesToCheck_13_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@12166.4]
  assign entriesToCheck_13_8 = _T_13242 & checkBits_13; // @[LoadQueue.scala 141:26:@12167.4]
  assign _T_13244 = storesToCheck_13_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@12168.4]
  assign entriesToCheck_13_9 = _T_13244 & checkBits_13; // @[LoadQueue.scala 141:26:@12169.4]
  assign _T_13246 = storesToCheck_13_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@12170.4]
  assign entriesToCheck_13_10 = _T_13246 & checkBits_13; // @[LoadQueue.scala 141:26:@12171.4]
  assign _T_13248 = storesToCheck_13_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@12172.4]
  assign entriesToCheck_13_11 = _T_13248 & checkBits_13; // @[LoadQueue.scala 141:26:@12173.4]
  assign _T_13250 = storesToCheck_13_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@12174.4]
  assign entriesToCheck_13_12 = _T_13250 & checkBits_13; // @[LoadQueue.scala 141:26:@12175.4]
  assign _T_13252 = storesToCheck_13_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@12176.4]
  assign entriesToCheck_13_13 = _T_13252 & checkBits_13; // @[LoadQueue.scala 141:26:@12177.4]
  assign _T_13254 = storesToCheck_13_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@12178.4]
  assign entriesToCheck_13_14 = _T_13254 & checkBits_13; // @[LoadQueue.scala 141:26:@12179.4]
  assign _T_13256 = storesToCheck_13_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@12180.4]
  assign entriesToCheck_13_15 = _T_13256 & checkBits_13; // @[LoadQueue.scala 141:26:@12181.4]
  assign _T_13258 = storesToCheck_14_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@12198.4]
  assign entriesToCheck_14_0 = _T_13258 & checkBits_14; // @[LoadQueue.scala 141:26:@12199.4]
  assign _T_13260 = storesToCheck_14_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@12200.4]
  assign entriesToCheck_14_1 = _T_13260 & checkBits_14; // @[LoadQueue.scala 141:26:@12201.4]
  assign _T_13262 = storesToCheck_14_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@12202.4]
  assign entriesToCheck_14_2 = _T_13262 & checkBits_14; // @[LoadQueue.scala 141:26:@12203.4]
  assign _T_13264 = storesToCheck_14_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@12204.4]
  assign entriesToCheck_14_3 = _T_13264 & checkBits_14; // @[LoadQueue.scala 141:26:@12205.4]
  assign _T_13266 = storesToCheck_14_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@12206.4]
  assign entriesToCheck_14_4 = _T_13266 & checkBits_14; // @[LoadQueue.scala 141:26:@12207.4]
  assign _T_13268 = storesToCheck_14_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@12208.4]
  assign entriesToCheck_14_5 = _T_13268 & checkBits_14; // @[LoadQueue.scala 141:26:@12209.4]
  assign _T_13270 = storesToCheck_14_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@12210.4]
  assign entriesToCheck_14_6 = _T_13270 & checkBits_14; // @[LoadQueue.scala 141:26:@12211.4]
  assign _T_13272 = storesToCheck_14_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@12212.4]
  assign entriesToCheck_14_7 = _T_13272 & checkBits_14; // @[LoadQueue.scala 141:26:@12213.4]
  assign _T_13274 = storesToCheck_14_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@12214.4]
  assign entriesToCheck_14_8 = _T_13274 & checkBits_14; // @[LoadQueue.scala 141:26:@12215.4]
  assign _T_13276 = storesToCheck_14_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@12216.4]
  assign entriesToCheck_14_9 = _T_13276 & checkBits_14; // @[LoadQueue.scala 141:26:@12217.4]
  assign _T_13278 = storesToCheck_14_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@12218.4]
  assign entriesToCheck_14_10 = _T_13278 & checkBits_14; // @[LoadQueue.scala 141:26:@12219.4]
  assign _T_13280 = storesToCheck_14_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@12220.4]
  assign entriesToCheck_14_11 = _T_13280 & checkBits_14; // @[LoadQueue.scala 141:26:@12221.4]
  assign _T_13282 = storesToCheck_14_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@12222.4]
  assign entriesToCheck_14_12 = _T_13282 & checkBits_14; // @[LoadQueue.scala 141:26:@12223.4]
  assign _T_13284 = storesToCheck_14_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@12224.4]
  assign entriesToCheck_14_13 = _T_13284 & checkBits_14; // @[LoadQueue.scala 141:26:@12225.4]
  assign _T_13286 = storesToCheck_14_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@12226.4]
  assign entriesToCheck_14_14 = _T_13286 & checkBits_14; // @[LoadQueue.scala 141:26:@12227.4]
  assign _T_13288 = storesToCheck_14_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@12228.4]
  assign entriesToCheck_14_15 = _T_13288 & checkBits_14; // @[LoadQueue.scala 141:26:@12229.4]
  assign _T_13290 = storesToCheck_15_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@12246.4]
  assign entriesToCheck_15_0 = _T_13290 & checkBits_15; // @[LoadQueue.scala 141:26:@12247.4]
  assign _T_13292 = storesToCheck_15_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@12248.4]
  assign entriesToCheck_15_1 = _T_13292 & checkBits_15; // @[LoadQueue.scala 141:26:@12249.4]
  assign _T_13294 = storesToCheck_15_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@12250.4]
  assign entriesToCheck_15_2 = _T_13294 & checkBits_15; // @[LoadQueue.scala 141:26:@12251.4]
  assign _T_13296 = storesToCheck_15_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@12252.4]
  assign entriesToCheck_15_3 = _T_13296 & checkBits_15; // @[LoadQueue.scala 141:26:@12253.4]
  assign _T_13298 = storesToCheck_15_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@12254.4]
  assign entriesToCheck_15_4 = _T_13298 & checkBits_15; // @[LoadQueue.scala 141:26:@12255.4]
  assign _T_13300 = storesToCheck_15_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@12256.4]
  assign entriesToCheck_15_5 = _T_13300 & checkBits_15; // @[LoadQueue.scala 141:26:@12257.4]
  assign _T_13302 = storesToCheck_15_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@12258.4]
  assign entriesToCheck_15_6 = _T_13302 & checkBits_15; // @[LoadQueue.scala 141:26:@12259.4]
  assign _T_13304 = storesToCheck_15_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@12260.4]
  assign entriesToCheck_15_7 = _T_13304 & checkBits_15; // @[LoadQueue.scala 141:26:@12261.4]
  assign _T_13306 = storesToCheck_15_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@12262.4]
  assign entriesToCheck_15_8 = _T_13306 & checkBits_15; // @[LoadQueue.scala 141:26:@12263.4]
  assign _T_13308 = storesToCheck_15_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@12264.4]
  assign entriesToCheck_15_9 = _T_13308 & checkBits_15; // @[LoadQueue.scala 141:26:@12265.4]
  assign _T_13310 = storesToCheck_15_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@12266.4]
  assign entriesToCheck_15_10 = _T_13310 & checkBits_15; // @[LoadQueue.scala 141:26:@12267.4]
  assign _T_13312 = storesToCheck_15_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@12268.4]
  assign entriesToCheck_15_11 = _T_13312 & checkBits_15; // @[LoadQueue.scala 141:26:@12269.4]
  assign _T_13314 = storesToCheck_15_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@12270.4]
  assign entriesToCheck_15_12 = _T_13314 & checkBits_15; // @[LoadQueue.scala 141:26:@12271.4]
  assign _T_13316 = storesToCheck_15_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@12272.4]
  assign entriesToCheck_15_13 = _T_13316 & checkBits_15; // @[LoadQueue.scala 141:26:@12273.4]
  assign _T_13318 = storesToCheck_15_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@12274.4]
  assign entriesToCheck_15_14 = _T_13318 & checkBits_15; // @[LoadQueue.scala 141:26:@12275.4]
  assign _T_13320 = storesToCheck_15_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@12276.4]
  assign entriesToCheck_15_15 = _T_13320 & checkBits_15; // @[LoadQueue.scala 141:26:@12277.4]
  assign _T_14552 = entriesToCheck_0_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12295.4]
  assign _T_14553 = _T_14552 & addrKnown_0; // @[LoadQueue.scala 152:41:@12296.4]
  assign _T_14554 = addrQ_0 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12297.4]
  assign conflict_0_0 = _T_14553 & _T_14554; // @[LoadQueue.scala 152:68:@12298.4]
  assign _T_14556 = entriesToCheck_0_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12300.4]
  assign _T_14557 = _T_14556 & addrKnown_0; // @[LoadQueue.scala 152:41:@12301.4]
  assign _T_14558 = addrQ_0 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12302.4]
  assign conflict_0_1 = _T_14557 & _T_14558; // @[LoadQueue.scala 152:68:@12303.4]
  assign _T_14560 = entriesToCheck_0_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12305.4]
  assign _T_14561 = _T_14560 & addrKnown_0; // @[LoadQueue.scala 152:41:@12306.4]
  assign _T_14562 = addrQ_0 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12307.4]
  assign conflict_0_2 = _T_14561 & _T_14562; // @[LoadQueue.scala 152:68:@12308.4]
  assign _T_14564 = entriesToCheck_0_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12310.4]
  assign _T_14565 = _T_14564 & addrKnown_0; // @[LoadQueue.scala 152:41:@12311.4]
  assign _T_14566 = addrQ_0 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12312.4]
  assign conflict_0_3 = _T_14565 & _T_14566; // @[LoadQueue.scala 152:68:@12313.4]
  assign _T_14568 = entriesToCheck_0_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12315.4]
  assign _T_14569 = _T_14568 & addrKnown_0; // @[LoadQueue.scala 152:41:@12316.4]
  assign _T_14570 = addrQ_0 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12317.4]
  assign conflict_0_4 = _T_14569 & _T_14570; // @[LoadQueue.scala 152:68:@12318.4]
  assign _T_14572 = entriesToCheck_0_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12320.4]
  assign _T_14573 = _T_14572 & addrKnown_0; // @[LoadQueue.scala 152:41:@12321.4]
  assign _T_14574 = addrQ_0 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12322.4]
  assign conflict_0_5 = _T_14573 & _T_14574; // @[LoadQueue.scala 152:68:@12323.4]
  assign _T_14576 = entriesToCheck_0_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12325.4]
  assign _T_14577 = _T_14576 & addrKnown_0; // @[LoadQueue.scala 152:41:@12326.4]
  assign _T_14578 = addrQ_0 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12327.4]
  assign conflict_0_6 = _T_14577 & _T_14578; // @[LoadQueue.scala 152:68:@12328.4]
  assign _T_14580 = entriesToCheck_0_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12330.4]
  assign _T_14581 = _T_14580 & addrKnown_0; // @[LoadQueue.scala 152:41:@12331.4]
  assign _T_14582 = addrQ_0 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12332.4]
  assign conflict_0_7 = _T_14581 & _T_14582; // @[LoadQueue.scala 152:68:@12333.4]
  assign _T_14584 = entriesToCheck_0_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12335.4]
  assign _T_14585 = _T_14584 & addrKnown_0; // @[LoadQueue.scala 152:41:@12336.4]
  assign _T_14586 = addrQ_0 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12337.4]
  assign conflict_0_8 = _T_14585 & _T_14586; // @[LoadQueue.scala 152:68:@12338.4]
  assign _T_14588 = entriesToCheck_0_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12340.4]
  assign _T_14589 = _T_14588 & addrKnown_0; // @[LoadQueue.scala 152:41:@12341.4]
  assign _T_14590 = addrQ_0 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12342.4]
  assign conflict_0_9 = _T_14589 & _T_14590; // @[LoadQueue.scala 152:68:@12343.4]
  assign _T_14592 = entriesToCheck_0_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12345.4]
  assign _T_14593 = _T_14592 & addrKnown_0; // @[LoadQueue.scala 152:41:@12346.4]
  assign _T_14594 = addrQ_0 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12347.4]
  assign conflict_0_10 = _T_14593 & _T_14594; // @[LoadQueue.scala 152:68:@12348.4]
  assign _T_14596 = entriesToCheck_0_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12350.4]
  assign _T_14597 = _T_14596 & addrKnown_0; // @[LoadQueue.scala 152:41:@12351.4]
  assign _T_14598 = addrQ_0 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12352.4]
  assign conflict_0_11 = _T_14597 & _T_14598; // @[LoadQueue.scala 152:68:@12353.4]
  assign _T_14600 = entriesToCheck_0_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12355.4]
  assign _T_14601 = _T_14600 & addrKnown_0; // @[LoadQueue.scala 152:41:@12356.4]
  assign _T_14602 = addrQ_0 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12357.4]
  assign conflict_0_12 = _T_14601 & _T_14602; // @[LoadQueue.scala 152:68:@12358.4]
  assign _T_14604 = entriesToCheck_0_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@12360.4]
  assign _T_14605 = _T_14604 & addrKnown_0; // @[LoadQueue.scala 152:41:@12361.4]
  assign _T_14606 = addrQ_0 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@12362.4]
  assign conflict_0_13 = _T_14605 & _T_14606; // @[LoadQueue.scala 152:68:@12363.4]
  assign _T_14608 = entriesToCheck_0_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@12365.4]
  assign _T_14609 = _T_14608 & addrKnown_0; // @[LoadQueue.scala 152:41:@12366.4]
  assign _T_14610 = addrQ_0 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@12367.4]
  assign conflict_0_14 = _T_14609 & _T_14610; // @[LoadQueue.scala 152:68:@12368.4]
  assign _T_14612 = entriesToCheck_0_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@12370.4]
  assign _T_14613 = _T_14612 & addrKnown_0; // @[LoadQueue.scala 152:41:@12371.4]
  assign _T_14614 = addrQ_0 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@12372.4]
  assign conflict_0_15 = _T_14613 & _T_14614; // @[LoadQueue.scala 152:68:@12373.4]
  assign _T_14616 = entriesToCheck_1_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12375.4]
  assign _T_14617 = _T_14616 & addrKnown_1; // @[LoadQueue.scala 152:41:@12376.4]
  assign _T_14618 = addrQ_1 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12377.4]
  assign conflict_1_0 = _T_14617 & _T_14618; // @[LoadQueue.scala 152:68:@12378.4]
  assign _T_14620 = entriesToCheck_1_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12380.4]
  assign _T_14621 = _T_14620 & addrKnown_1; // @[LoadQueue.scala 152:41:@12381.4]
  assign _T_14622 = addrQ_1 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12382.4]
  assign conflict_1_1 = _T_14621 & _T_14622; // @[LoadQueue.scala 152:68:@12383.4]
  assign _T_14624 = entriesToCheck_1_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12385.4]
  assign _T_14625 = _T_14624 & addrKnown_1; // @[LoadQueue.scala 152:41:@12386.4]
  assign _T_14626 = addrQ_1 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12387.4]
  assign conflict_1_2 = _T_14625 & _T_14626; // @[LoadQueue.scala 152:68:@12388.4]
  assign _T_14628 = entriesToCheck_1_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12390.4]
  assign _T_14629 = _T_14628 & addrKnown_1; // @[LoadQueue.scala 152:41:@12391.4]
  assign _T_14630 = addrQ_1 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12392.4]
  assign conflict_1_3 = _T_14629 & _T_14630; // @[LoadQueue.scala 152:68:@12393.4]
  assign _T_14632 = entriesToCheck_1_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12395.4]
  assign _T_14633 = _T_14632 & addrKnown_1; // @[LoadQueue.scala 152:41:@12396.4]
  assign _T_14634 = addrQ_1 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12397.4]
  assign conflict_1_4 = _T_14633 & _T_14634; // @[LoadQueue.scala 152:68:@12398.4]
  assign _T_14636 = entriesToCheck_1_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12400.4]
  assign _T_14637 = _T_14636 & addrKnown_1; // @[LoadQueue.scala 152:41:@12401.4]
  assign _T_14638 = addrQ_1 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12402.4]
  assign conflict_1_5 = _T_14637 & _T_14638; // @[LoadQueue.scala 152:68:@12403.4]
  assign _T_14640 = entriesToCheck_1_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12405.4]
  assign _T_14641 = _T_14640 & addrKnown_1; // @[LoadQueue.scala 152:41:@12406.4]
  assign _T_14642 = addrQ_1 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12407.4]
  assign conflict_1_6 = _T_14641 & _T_14642; // @[LoadQueue.scala 152:68:@12408.4]
  assign _T_14644 = entriesToCheck_1_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12410.4]
  assign _T_14645 = _T_14644 & addrKnown_1; // @[LoadQueue.scala 152:41:@12411.4]
  assign _T_14646 = addrQ_1 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12412.4]
  assign conflict_1_7 = _T_14645 & _T_14646; // @[LoadQueue.scala 152:68:@12413.4]
  assign _T_14648 = entriesToCheck_1_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12415.4]
  assign _T_14649 = _T_14648 & addrKnown_1; // @[LoadQueue.scala 152:41:@12416.4]
  assign _T_14650 = addrQ_1 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12417.4]
  assign conflict_1_8 = _T_14649 & _T_14650; // @[LoadQueue.scala 152:68:@12418.4]
  assign _T_14652 = entriesToCheck_1_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12420.4]
  assign _T_14653 = _T_14652 & addrKnown_1; // @[LoadQueue.scala 152:41:@12421.4]
  assign _T_14654 = addrQ_1 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12422.4]
  assign conflict_1_9 = _T_14653 & _T_14654; // @[LoadQueue.scala 152:68:@12423.4]
  assign _T_14656 = entriesToCheck_1_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12425.4]
  assign _T_14657 = _T_14656 & addrKnown_1; // @[LoadQueue.scala 152:41:@12426.4]
  assign _T_14658 = addrQ_1 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12427.4]
  assign conflict_1_10 = _T_14657 & _T_14658; // @[LoadQueue.scala 152:68:@12428.4]
  assign _T_14660 = entriesToCheck_1_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12430.4]
  assign _T_14661 = _T_14660 & addrKnown_1; // @[LoadQueue.scala 152:41:@12431.4]
  assign _T_14662 = addrQ_1 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12432.4]
  assign conflict_1_11 = _T_14661 & _T_14662; // @[LoadQueue.scala 152:68:@12433.4]
  assign _T_14664 = entriesToCheck_1_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12435.4]
  assign _T_14665 = _T_14664 & addrKnown_1; // @[LoadQueue.scala 152:41:@12436.4]
  assign _T_14666 = addrQ_1 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12437.4]
  assign conflict_1_12 = _T_14665 & _T_14666; // @[LoadQueue.scala 152:68:@12438.4]
  assign _T_14668 = entriesToCheck_1_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@12440.4]
  assign _T_14669 = _T_14668 & addrKnown_1; // @[LoadQueue.scala 152:41:@12441.4]
  assign _T_14670 = addrQ_1 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@12442.4]
  assign conflict_1_13 = _T_14669 & _T_14670; // @[LoadQueue.scala 152:68:@12443.4]
  assign _T_14672 = entriesToCheck_1_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@12445.4]
  assign _T_14673 = _T_14672 & addrKnown_1; // @[LoadQueue.scala 152:41:@12446.4]
  assign _T_14674 = addrQ_1 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@12447.4]
  assign conflict_1_14 = _T_14673 & _T_14674; // @[LoadQueue.scala 152:68:@12448.4]
  assign _T_14676 = entriesToCheck_1_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@12450.4]
  assign _T_14677 = _T_14676 & addrKnown_1; // @[LoadQueue.scala 152:41:@12451.4]
  assign _T_14678 = addrQ_1 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@12452.4]
  assign conflict_1_15 = _T_14677 & _T_14678; // @[LoadQueue.scala 152:68:@12453.4]
  assign _T_14680 = entriesToCheck_2_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12455.4]
  assign _T_14681 = _T_14680 & addrKnown_2; // @[LoadQueue.scala 152:41:@12456.4]
  assign _T_14682 = addrQ_2 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12457.4]
  assign conflict_2_0 = _T_14681 & _T_14682; // @[LoadQueue.scala 152:68:@12458.4]
  assign _T_14684 = entriesToCheck_2_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12460.4]
  assign _T_14685 = _T_14684 & addrKnown_2; // @[LoadQueue.scala 152:41:@12461.4]
  assign _T_14686 = addrQ_2 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12462.4]
  assign conflict_2_1 = _T_14685 & _T_14686; // @[LoadQueue.scala 152:68:@12463.4]
  assign _T_14688 = entriesToCheck_2_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12465.4]
  assign _T_14689 = _T_14688 & addrKnown_2; // @[LoadQueue.scala 152:41:@12466.4]
  assign _T_14690 = addrQ_2 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12467.4]
  assign conflict_2_2 = _T_14689 & _T_14690; // @[LoadQueue.scala 152:68:@12468.4]
  assign _T_14692 = entriesToCheck_2_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12470.4]
  assign _T_14693 = _T_14692 & addrKnown_2; // @[LoadQueue.scala 152:41:@12471.4]
  assign _T_14694 = addrQ_2 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12472.4]
  assign conflict_2_3 = _T_14693 & _T_14694; // @[LoadQueue.scala 152:68:@12473.4]
  assign _T_14696 = entriesToCheck_2_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12475.4]
  assign _T_14697 = _T_14696 & addrKnown_2; // @[LoadQueue.scala 152:41:@12476.4]
  assign _T_14698 = addrQ_2 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12477.4]
  assign conflict_2_4 = _T_14697 & _T_14698; // @[LoadQueue.scala 152:68:@12478.4]
  assign _T_14700 = entriesToCheck_2_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12480.4]
  assign _T_14701 = _T_14700 & addrKnown_2; // @[LoadQueue.scala 152:41:@12481.4]
  assign _T_14702 = addrQ_2 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12482.4]
  assign conflict_2_5 = _T_14701 & _T_14702; // @[LoadQueue.scala 152:68:@12483.4]
  assign _T_14704 = entriesToCheck_2_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12485.4]
  assign _T_14705 = _T_14704 & addrKnown_2; // @[LoadQueue.scala 152:41:@12486.4]
  assign _T_14706 = addrQ_2 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12487.4]
  assign conflict_2_6 = _T_14705 & _T_14706; // @[LoadQueue.scala 152:68:@12488.4]
  assign _T_14708 = entriesToCheck_2_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12490.4]
  assign _T_14709 = _T_14708 & addrKnown_2; // @[LoadQueue.scala 152:41:@12491.4]
  assign _T_14710 = addrQ_2 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12492.4]
  assign conflict_2_7 = _T_14709 & _T_14710; // @[LoadQueue.scala 152:68:@12493.4]
  assign _T_14712 = entriesToCheck_2_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12495.4]
  assign _T_14713 = _T_14712 & addrKnown_2; // @[LoadQueue.scala 152:41:@12496.4]
  assign _T_14714 = addrQ_2 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12497.4]
  assign conflict_2_8 = _T_14713 & _T_14714; // @[LoadQueue.scala 152:68:@12498.4]
  assign _T_14716 = entriesToCheck_2_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12500.4]
  assign _T_14717 = _T_14716 & addrKnown_2; // @[LoadQueue.scala 152:41:@12501.4]
  assign _T_14718 = addrQ_2 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12502.4]
  assign conflict_2_9 = _T_14717 & _T_14718; // @[LoadQueue.scala 152:68:@12503.4]
  assign _T_14720 = entriesToCheck_2_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12505.4]
  assign _T_14721 = _T_14720 & addrKnown_2; // @[LoadQueue.scala 152:41:@12506.4]
  assign _T_14722 = addrQ_2 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12507.4]
  assign conflict_2_10 = _T_14721 & _T_14722; // @[LoadQueue.scala 152:68:@12508.4]
  assign _T_14724 = entriesToCheck_2_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12510.4]
  assign _T_14725 = _T_14724 & addrKnown_2; // @[LoadQueue.scala 152:41:@12511.4]
  assign _T_14726 = addrQ_2 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12512.4]
  assign conflict_2_11 = _T_14725 & _T_14726; // @[LoadQueue.scala 152:68:@12513.4]
  assign _T_14728 = entriesToCheck_2_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12515.4]
  assign _T_14729 = _T_14728 & addrKnown_2; // @[LoadQueue.scala 152:41:@12516.4]
  assign _T_14730 = addrQ_2 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12517.4]
  assign conflict_2_12 = _T_14729 & _T_14730; // @[LoadQueue.scala 152:68:@12518.4]
  assign _T_14732 = entriesToCheck_2_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@12520.4]
  assign _T_14733 = _T_14732 & addrKnown_2; // @[LoadQueue.scala 152:41:@12521.4]
  assign _T_14734 = addrQ_2 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@12522.4]
  assign conflict_2_13 = _T_14733 & _T_14734; // @[LoadQueue.scala 152:68:@12523.4]
  assign _T_14736 = entriesToCheck_2_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@12525.4]
  assign _T_14737 = _T_14736 & addrKnown_2; // @[LoadQueue.scala 152:41:@12526.4]
  assign _T_14738 = addrQ_2 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@12527.4]
  assign conflict_2_14 = _T_14737 & _T_14738; // @[LoadQueue.scala 152:68:@12528.4]
  assign _T_14740 = entriesToCheck_2_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@12530.4]
  assign _T_14741 = _T_14740 & addrKnown_2; // @[LoadQueue.scala 152:41:@12531.4]
  assign _T_14742 = addrQ_2 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@12532.4]
  assign conflict_2_15 = _T_14741 & _T_14742; // @[LoadQueue.scala 152:68:@12533.4]
  assign _T_14744 = entriesToCheck_3_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12535.4]
  assign _T_14745 = _T_14744 & addrKnown_3; // @[LoadQueue.scala 152:41:@12536.4]
  assign _T_14746 = addrQ_3 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12537.4]
  assign conflict_3_0 = _T_14745 & _T_14746; // @[LoadQueue.scala 152:68:@12538.4]
  assign _T_14748 = entriesToCheck_3_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12540.4]
  assign _T_14749 = _T_14748 & addrKnown_3; // @[LoadQueue.scala 152:41:@12541.4]
  assign _T_14750 = addrQ_3 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12542.4]
  assign conflict_3_1 = _T_14749 & _T_14750; // @[LoadQueue.scala 152:68:@12543.4]
  assign _T_14752 = entriesToCheck_3_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12545.4]
  assign _T_14753 = _T_14752 & addrKnown_3; // @[LoadQueue.scala 152:41:@12546.4]
  assign _T_14754 = addrQ_3 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12547.4]
  assign conflict_3_2 = _T_14753 & _T_14754; // @[LoadQueue.scala 152:68:@12548.4]
  assign _T_14756 = entriesToCheck_3_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12550.4]
  assign _T_14757 = _T_14756 & addrKnown_3; // @[LoadQueue.scala 152:41:@12551.4]
  assign _T_14758 = addrQ_3 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12552.4]
  assign conflict_3_3 = _T_14757 & _T_14758; // @[LoadQueue.scala 152:68:@12553.4]
  assign _T_14760 = entriesToCheck_3_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12555.4]
  assign _T_14761 = _T_14760 & addrKnown_3; // @[LoadQueue.scala 152:41:@12556.4]
  assign _T_14762 = addrQ_3 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12557.4]
  assign conflict_3_4 = _T_14761 & _T_14762; // @[LoadQueue.scala 152:68:@12558.4]
  assign _T_14764 = entriesToCheck_3_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12560.4]
  assign _T_14765 = _T_14764 & addrKnown_3; // @[LoadQueue.scala 152:41:@12561.4]
  assign _T_14766 = addrQ_3 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12562.4]
  assign conflict_3_5 = _T_14765 & _T_14766; // @[LoadQueue.scala 152:68:@12563.4]
  assign _T_14768 = entriesToCheck_3_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12565.4]
  assign _T_14769 = _T_14768 & addrKnown_3; // @[LoadQueue.scala 152:41:@12566.4]
  assign _T_14770 = addrQ_3 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12567.4]
  assign conflict_3_6 = _T_14769 & _T_14770; // @[LoadQueue.scala 152:68:@12568.4]
  assign _T_14772 = entriesToCheck_3_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12570.4]
  assign _T_14773 = _T_14772 & addrKnown_3; // @[LoadQueue.scala 152:41:@12571.4]
  assign _T_14774 = addrQ_3 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12572.4]
  assign conflict_3_7 = _T_14773 & _T_14774; // @[LoadQueue.scala 152:68:@12573.4]
  assign _T_14776 = entriesToCheck_3_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12575.4]
  assign _T_14777 = _T_14776 & addrKnown_3; // @[LoadQueue.scala 152:41:@12576.4]
  assign _T_14778 = addrQ_3 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12577.4]
  assign conflict_3_8 = _T_14777 & _T_14778; // @[LoadQueue.scala 152:68:@12578.4]
  assign _T_14780 = entriesToCheck_3_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12580.4]
  assign _T_14781 = _T_14780 & addrKnown_3; // @[LoadQueue.scala 152:41:@12581.4]
  assign _T_14782 = addrQ_3 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12582.4]
  assign conflict_3_9 = _T_14781 & _T_14782; // @[LoadQueue.scala 152:68:@12583.4]
  assign _T_14784 = entriesToCheck_3_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12585.4]
  assign _T_14785 = _T_14784 & addrKnown_3; // @[LoadQueue.scala 152:41:@12586.4]
  assign _T_14786 = addrQ_3 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12587.4]
  assign conflict_3_10 = _T_14785 & _T_14786; // @[LoadQueue.scala 152:68:@12588.4]
  assign _T_14788 = entriesToCheck_3_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12590.4]
  assign _T_14789 = _T_14788 & addrKnown_3; // @[LoadQueue.scala 152:41:@12591.4]
  assign _T_14790 = addrQ_3 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12592.4]
  assign conflict_3_11 = _T_14789 & _T_14790; // @[LoadQueue.scala 152:68:@12593.4]
  assign _T_14792 = entriesToCheck_3_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12595.4]
  assign _T_14793 = _T_14792 & addrKnown_3; // @[LoadQueue.scala 152:41:@12596.4]
  assign _T_14794 = addrQ_3 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12597.4]
  assign conflict_3_12 = _T_14793 & _T_14794; // @[LoadQueue.scala 152:68:@12598.4]
  assign _T_14796 = entriesToCheck_3_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@12600.4]
  assign _T_14797 = _T_14796 & addrKnown_3; // @[LoadQueue.scala 152:41:@12601.4]
  assign _T_14798 = addrQ_3 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@12602.4]
  assign conflict_3_13 = _T_14797 & _T_14798; // @[LoadQueue.scala 152:68:@12603.4]
  assign _T_14800 = entriesToCheck_3_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@12605.4]
  assign _T_14801 = _T_14800 & addrKnown_3; // @[LoadQueue.scala 152:41:@12606.4]
  assign _T_14802 = addrQ_3 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@12607.4]
  assign conflict_3_14 = _T_14801 & _T_14802; // @[LoadQueue.scala 152:68:@12608.4]
  assign _T_14804 = entriesToCheck_3_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@12610.4]
  assign _T_14805 = _T_14804 & addrKnown_3; // @[LoadQueue.scala 152:41:@12611.4]
  assign _T_14806 = addrQ_3 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@12612.4]
  assign conflict_3_15 = _T_14805 & _T_14806; // @[LoadQueue.scala 152:68:@12613.4]
  assign _T_14808 = entriesToCheck_4_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12615.4]
  assign _T_14809 = _T_14808 & addrKnown_4; // @[LoadQueue.scala 152:41:@12616.4]
  assign _T_14810 = addrQ_4 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12617.4]
  assign conflict_4_0 = _T_14809 & _T_14810; // @[LoadQueue.scala 152:68:@12618.4]
  assign _T_14812 = entriesToCheck_4_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12620.4]
  assign _T_14813 = _T_14812 & addrKnown_4; // @[LoadQueue.scala 152:41:@12621.4]
  assign _T_14814 = addrQ_4 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12622.4]
  assign conflict_4_1 = _T_14813 & _T_14814; // @[LoadQueue.scala 152:68:@12623.4]
  assign _T_14816 = entriesToCheck_4_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12625.4]
  assign _T_14817 = _T_14816 & addrKnown_4; // @[LoadQueue.scala 152:41:@12626.4]
  assign _T_14818 = addrQ_4 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12627.4]
  assign conflict_4_2 = _T_14817 & _T_14818; // @[LoadQueue.scala 152:68:@12628.4]
  assign _T_14820 = entriesToCheck_4_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12630.4]
  assign _T_14821 = _T_14820 & addrKnown_4; // @[LoadQueue.scala 152:41:@12631.4]
  assign _T_14822 = addrQ_4 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12632.4]
  assign conflict_4_3 = _T_14821 & _T_14822; // @[LoadQueue.scala 152:68:@12633.4]
  assign _T_14824 = entriesToCheck_4_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12635.4]
  assign _T_14825 = _T_14824 & addrKnown_4; // @[LoadQueue.scala 152:41:@12636.4]
  assign _T_14826 = addrQ_4 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12637.4]
  assign conflict_4_4 = _T_14825 & _T_14826; // @[LoadQueue.scala 152:68:@12638.4]
  assign _T_14828 = entriesToCheck_4_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12640.4]
  assign _T_14829 = _T_14828 & addrKnown_4; // @[LoadQueue.scala 152:41:@12641.4]
  assign _T_14830 = addrQ_4 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12642.4]
  assign conflict_4_5 = _T_14829 & _T_14830; // @[LoadQueue.scala 152:68:@12643.4]
  assign _T_14832 = entriesToCheck_4_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12645.4]
  assign _T_14833 = _T_14832 & addrKnown_4; // @[LoadQueue.scala 152:41:@12646.4]
  assign _T_14834 = addrQ_4 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12647.4]
  assign conflict_4_6 = _T_14833 & _T_14834; // @[LoadQueue.scala 152:68:@12648.4]
  assign _T_14836 = entriesToCheck_4_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12650.4]
  assign _T_14837 = _T_14836 & addrKnown_4; // @[LoadQueue.scala 152:41:@12651.4]
  assign _T_14838 = addrQ_4 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12652.4]
  assign conflict_4_7 = _T_14837 & _T_14838; // @[LoadQueue.scala 152:68:@12653.4]
  assign _T_14840 = entriesToCheck_4_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12655.4]
  assign _T_14841 = _T_14840 & addrKnown_4; // @[LoadQueue.scala 152:41:@12656.4]
  assign _T_14842 = addrQ_4 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12657.4]
  assign conflict_4_8 = _T_14841 & _T_14842; // @[LoadQueue.scala 152:68:@12658.4]
  assign _T_14844 = entriesToCheck_4_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12660.4]
  assign _T_14845 = _T_14844 & addrKnown_4; // @[LoadQueue.scala 152:41:@12661.4]
  assign _T_14846 = addrQ_4 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12662.4]
  assign conflict_4_9 = _T_14845 & _T_14846; // @[LoadQueue.scala 152:68:@12663.4]
  assign _T_14848 = entriesToCheck_4_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12665.4]
  assign _T_14849 = _T_14848 & addrKnown_4; // @[LoadQueue.scala 152:41:@12666.4]
  assign _T_14850 = addrQ_4 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12667.4]
  assign conflict_4_10 = _T_14849 & _T_14850; // @[LoadQueue.scala 152:68:@12668.4]
  assign _T_14852 = entriesToCheck_4_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12670.4]
  assign _T_14853 = _T_14852 & addrKnown_4; // @[LoadQueue.scala 152:41:@12671.4]
  assign _T_14854 = addrQ_4 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12672.4]
  assign conflict_4_11 = _T_14853 & _T_14854; // @[LoadQueue.scala 152:68:@12673.4]
  assign _T_14856 = entriesToCheck_4_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12675.4]
  assign _T_14857 = _T_14856 & addrKnown_4; // @[LoadQueue.scala 152:41:@12676.4]
  assign _T_14858 = addrQ_4 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12677.4]
  assign conflict_4_12 = _T_14857 & _T_14858; // @[LoadQueue.scala 152:68:@12678.4]
  assign _T_14860 = entriesToCheck_4_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@12680.4]
  assign _T_14861 = _T_14860 & addrKnown_4; // @[LoadQueue.scala 152:41:@12681.4]
  assign _T_14862 = addrQ_4 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@12682.4]
  assign conflict_4_13 = _T_14861 & _T_14862; // @[LoadQueue.scala 152:68:@12683.4]
  assign _T_14864 = entriesToCheck_4_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@12685.4]
  assign _T_14865 = _T_14864 & addrKnown_4; // @[LoadQueue.scala 152:41:@12686.4]
  assign _T_14866 = addrQ_4 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@12687.4]
  assign conflict_4_14 = _T_14865 & _T_14866; // @[LoadQueue.scala 152:68:@12688.4]
  assign _T_14868 = entriesToCheck_4_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@12690.4]
  assign _T_14869 = _T_14868 & addrKnown_4; // @[LoadQueue.scala 152:41:@12691.4]
  assign _T_14870 = addrQ_4 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@12692.4]
  assign conflict_4_15 = _T_14869 & _T_14870; // @[LoadQueue.scala 152:68:@12693.4]
  assign _T_14872 = entriesToCheck_5_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12695.4]
  assign _T_14873 = _T_14872 & addrKnown_5; // @[LoadQueue.scala 152:41:@12696.4]
  assign _T_14874 = addrQ_5 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12697.4]
  assign conflict_5_0 = _T_14873 & _T_14874; // @[LoadQueue.scala 152:68:@12698.4]
  assign _T_14876 = entriesToCheck_5_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12700.4]
  assign _T_14877 = _T_14876 & addrKnown_5; // @[LoadQueue.scala 152:41:@12701.4]
  assign _T_14878 = addrQ_5 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12702.4]
  assign conflict_5_1 = _T_14877 & _T_14878; // @[LoadQueue.scala 152:68:@12703.4]
  assign _T_14880 = entriesToCheck_5_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12705.4]
  assign _T_14881 = _T_14880 & addrKnown_5; // @[LoadQueue.scala 152:41:@12706.4]
  assign _T_14882 = addrQ_5 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12707.4]
  assign conflict_5_2 = _T_14881 & _T_14882; // @[LoadQueue.scala 152:68:@12708.4]
  assign _T_14884 = entriesToCheck_5_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12710.4]
  assign _T_14885 = _T_14884 & addrKnown_5; // @[LoadQueue.scala 152:41:@12711.4]
  assign _T_14886 = addrQ_5 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12712.4]
  assign conflict_5_3 = _T_14885 & _T_14886; // @[LoadQueue.scala 152:68:@12713.4]
  assign _T_14888 = entriesToCheck_5_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12715.4]
  assign _T_14889 = _T_14888 & addrKnown_5; // @[LoadQueue.scala 152:41:@12716.4]
  assign _T_14890 = addrQ_5 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12717.4]
  assign conflict_5_4 = _T_14889 & _T_14890; // @[LoadQueue.scala 152:68:@12718.4]
  assign _T_14892 = entriesToCheck_5_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12720.4]
  assign _T_14893 = _T_14892 & addrKnown_5; // @[LoadQueue.scala 152:41:@12721.4]
  assign _T_14894 = addrQ_5 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12722.4]
  assign conflict_5_5 = _T_14893 & _T_14894; // @[LoadQueue.scala 152:68:@12723.4]
  assign _T_14896 = entriesToCheck_5_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12725.4]
  assign _T_14897 = _T_14896 & addrKnown_5; // @[LoadQueue.scala 152:41:@12726.4]
  assign _T_14898 = addrQ_5 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12727.4]
  assign conflict_5_6 = _T_14897 & _T_14898; // @[LoadQueue.scala 152:68:@12728.4]
  assign _T_14900 = entriesToCheck_5_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12730.4]
  assign _T_14901 = _T_14900 & addrKnown_5; // @[LoadQueue.scala 152:41:@12731.4]
  assign _T_14902 = addrQ_5 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12732.4]
  assign conflict_5_7 = _T_14901 & _T_14902; // @[LoadQueue.scala 152:68:@12733.4]
  assign _T_14904 = entriesToCheck_5_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12735.4]
  assign _T_14905 = _T_14904 & addrKnown_5; // @[LoadQueue.scala 152:41:@12736.4]
  assign _T_14906 = addrQ_5 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12737.4]
  assign conflict_5_8 = _T_14905 & _T_14906; // @[LoadQueue.scala 152:68:@12738.4]
  assign _T_14908 = entriesToCheck_5_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12740.4]
  assign _T_14909 = _T_14908 & addrKnown_5; // @[LoadQueue.scala 152:41:@12741.4]
  assign _T_14910 = addrQ_5 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12742.4]
  assign conflict_5_9 = _T_14909 & _T_14910; // @[LoadQueue.scala 152:68:@12743.4]
  assign _T_14912 = entriesToCheck_5_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12745.4]
  assign _T_14913 = _T_14912 & addrKnown_5; // @[LoadQueue.scala 152:41:@12746.4]
  assign _T_14914 = addrQ_5 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12747.4]
  assign conflict_5_10 = _T_14913 & _T_14914; // @[LoadQueue.scala 152:68:@12748.4]
  assign _T_14916 = entriesToCheck_5_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12750.4]
  assign _T_14917 = _T_14916 & addrKnown_5; // @[LoadQueue.scala 152:41:@12751.4]
  assign _T_14918 = addrQ_5 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12752.4]
  assign conflict_5_11 = _T_14917 & _T_14918; // @[LoadQueue.scala 152:68:@12753.4]
  assign _T_14920 = entriesToCheck_5_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12755.4]
  assign _T_14921 = _T_14920 & addrKnown_5; // @[LoadQueue.scala 152:41:@12756.4]
  assign _T_14922 = addrQ_5 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12757.4]
  assign conflict_5_12 = _T_14921 & _T_14922; // @[LoadQueue.scala 152:68:@12758.4]
  assign _T_14924 = entriesToCheck_5_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@12760.4]
  assign _T_14925 = _T_14924 & addrKnown_5; // @[LoadQueue.scala 152:41:@12761.4]
  assign _T_14926 = addrQ_5 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@12762.4]
  assign conflict_5_13 = _T_14925 & _T_14926; // @[LoadQueue.scala 152:68:@12763.4]
  assign _T_14928 = entriesToCheck_5_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@12765.4]
  assign _T_14929 = _T_14928 & addrKnown_5; // @[LoadQueue.scala 152:41:@12766.4]
  assign _T_14930 = addrQ_5 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@12767.4]
  assign conflict_5_14 = _T_14929 & _T_14930; // @[LoadQueue.scala 152:68:@12768.4]
  assign _T_14932 = entriesToCheck_5_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@12770.4]
  assign _T_14933 = _T_14932 & addrKnown_5; // @[LoadQueue.scala 152:41:@12771.4]
  assign _T_14934 = addrQ_5 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@12772.4]
  assign conflict_5_15 = _T_14933 & _T_14934; // @[LoadQueue.scala 152:68:@12773.4]
  assign _T_14936 = entriesToCheck_6_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12775.4]
  assign _T_14937 = _T_14936 & addrKnown_6; // @[LoadQueue.scala 152:41:@12776.4]
  assign _T_14938 = addrQ_6 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12777.4]
  assign conflict_6_0 = _T_14937 & _T_14938; // @[LoadQueue.scala 152:68:@12778.4]
  assign _T_14940 = entriesToCheck_6_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12780.4]
  assign _T_14941 = _T_14940 & addrKnown_6; // @[LoadQueue.scala 152:41:@12781.4]
  assign _T_14942 = addrQ_6 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12782.4]
  assign conflict_6_1 = _T_14941 & _T_14942; // @[LoadQueue.scala 152:68:@12783.4]
  assign _T_14944 = entriesToCheck_6_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12785.4]
  assign _T_14945 = _T_14944 & addrKnown_6; // @[LoadQueue.scala 152:41:@12786.4]
  assign _T_14946 = addrQ_6 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12787.4]
  assign conflict_6_2 = _T_14945 & _T_14946; // @[LoadQueue.scala 152:68:@12788.4]
  assign _T_14948 = entriesToCheck_6_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12790.4]
  assign _T_14949 = _T_14948 & addrKnown_6; // @[LoadQueue.scala 152:41:@12791.4]
  assign _T_14950 = addrQ_6 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12792.4]
  assign conflict_6_3 = _T_14949 & _T_14950; // @[LoadQueue.scala 152:68:@12793.4]
  assign _T_14952 = entriesToCheck_6_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12795.4]
  assign _T_14953 = _T_14952 & addrKnown_6; // @[LoadQueue.scala 152:41:@12796.4]
  assign _T_14954 = addrQ_6 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12797.4]
  assign conflict_6_4 = _T_14953 & _T_14954; // @[LoadQueue.scala 152:68:@12798.4]
  assign _T_14956 = entriesToCheck_6_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12800.4]
  assign _T_14957 = _T_14956 & addrKnown_6; // @[LoadQueue.scala 152:41:@12801.4]
  assign _T_14958 = addrQ_6 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12802.4]
  assign conflict_6_5 = _T_14957 & _T_14958; // @[LoadQueue.scala 152:68:@12803.4]
  assign _T_14960 = entriesToCheck_6_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12805.4]
  assign _T_14961 = _T_14960 & addrKnown_6; // @[LoadQueue.scala 152:41:@12806.4]
  assign _T_14962 = addrQ_6 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12807.4]
  assign conflict_6_6 = _T_14961 & _T_14962; // @[LoadQueue.scala 152:68:@12808.4]
  assign _T_14964 = entriesToCheck_6_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12810.4]
  assign _T_14965 = _T_14964 & addrKnown_6; // @[LoadQueue.scala 152:41:@12811.4]
  assign _T_14966 = addrQ_6 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12812.4]
  assign conflict_6_7 = _T_14965 & _T_14966; // @[LoadQueue.scala 152:68:@12813.4]
  assign _T_14968 = entriesToCheck_6_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12815.4]
  assign _T_14969 = _T_14968 & addrKnown_6; // @[LoadQueue.scala 152:41:@12816.4]
  assign _T_14970 = addrQ_6 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12817.4]
  assign conflict_6_8 = _T_14969 & _T_14970; // @[LoadQueue.scala 152:68:@12818.4]
  assign _T_14972 = entriesToCheck_6_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12820.4]
  assign _T_14973 = _T_14972 & addrKnown_6; // @[LoadQueue.scala 152:41:@12821.4]
  assign _T_14974 = addrQ_6 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12822.4]
  assign conflict_6_9 = _T_14973 & _T_14974; // @[LoadQueue.scala 152:68:@12823.4]
  assign _T_14976 = entriesToCheck_6_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12825.4]
  assign _T_14977 = _T_14976 & addrKnown_6; // @[LoadQueue.scala 152:41:@12826.4]
  assign _T_14978 = addrQ_6 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12827.4]
  assign conflict_6_10 = _T_14977 & _T_14978; // @[LoadQueue.scala 152:68:@12828.4]
  assign _T_14980 = entriesToCheck_6_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12830.4]
  assign _T_14981 = _T_14980 & addrKnown_6; // @[LoadQueue.scala 152:41:@12831.4]
  assign _T_14982 = addrQ_6 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12832.4]
  assign conflict_6_11 = _T_14981 & _T_14982; // @[LoadQueue.scala 152:68:@12833.4]
  assign _T_14984 = entriesToCheck_6_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12835.4]
  assign _T_14985 = _T_14984 & addrKnown_6; // @[LoadQueue.scala 152:41:@12836.4]
  assign _T_14986 = addrQ_6 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12837.4]
  assign conflict_6_12 = _T_14985 & _T_14986; // @[LoadQueue.scala 152:68:@12838.4]
  assign _T_14988 = entriesToCheck_6_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@12840.4]
  assign _T_14989 = _T_14988 & addrKnown_6; // @[LoadQueue.scala 152:41:@12841.4]
  assign _T_14990 = addrQ_6 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@12842.4]
  assign conflict_6_13 = _T_14989 & _T_14990; // @[LoadQueue.scala 152:68:@12843.4]
  assign _T_14992 = entriesToCheck_6_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@12845.4]
  assign _T_14993 = _T_14992 & addrKnown_6; // @[LoadQueue.scala 152:41:@12846.4]
  assign _T_14994 = addrQ_6 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@12847.4]
  assign conflict_6_14 = _T_14993 & _T_14994; // @[LoadQueue.scala 152:68:@12848.4]
  assign _T_14996 = entriesToCheck_6_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@12850.4]
  assign _T_14997 = _T_14996 & addrKnown_6; // @[LoadQueue.scala 152:41:@12851.4]
  assign _T_14998 = addrQ_6 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@12852.4]
  assign conflict_6_15 = _T_14997 & _T_14998; // @[LoadQueue.scala 152:68:@12853.4]
  assign _T_15000 = entriesToCheck_7_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12855.4]
  assign _T_15001 = _T_15000 & addrKnown_7; // @[LoadQueue.scala 152:41:@12856.4]
  assign _T_15002 = addrQ_7 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12857.4]
  assign conflict_7_0 = _T_15001 & _T_15002; // @[LoadQueue.scala 152:68:@12858.4]
  assign _T_15004 = entriesToCheck_7_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12860.4]
  assign _T_15005 = _T_15004 & addrKnown_7; // @[LoadQueue.scala 152:41:@12861.4]
  assign _T_15006 = addrQ_7 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12862.4]
  assign conflict_7_1 = _T_15005 & _T_15006; // @[LoadQueue.scala 152:68:@12863.4]
  assign _T_15008 = entriesToCheck_7_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12865.4]
  assign _T_15009 = _T_15008 & addrKnown_7; // @[LoadQueue.scala 152:41:@12866.4]
  assign _T_15010 = addrQ_7 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12867.4]
  assign conflict_7_2 = _T_15009 & _T_15010; // @[LoadQueue.scala 152:68:@12868.4]
  assign _T_15012 = entriesToCheck_7_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12870.4]
  assign _T_15013 = _T_15012 & addrKnown_7; // @[LoadQueue.scala 152:41:@12871.4]
  assign _T_15014 = addrQ_7 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12872.4]
  assign conflict_7_3 = _T_15013 & _T_15014; // @[LoadQueue.scala 152:68:@12873.4]
  assign _T_15016 = entriesToCheck_7_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12875.4]
  assign _T_15017 = _T_15016 & addrKnown_7; // @[LoadQueue.scala 152:41:@12876.4]
  assign _T_15018 = addrQ_7 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12877.4]
  assign conflict_7_4 = _T_15017 & _T_15018; // @[LoadQueue.scala 152:68:@12878.4]
  assign _T_15020 = entriesToCheck_7_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12880.4]
  assign _T_15021 = _T_15020 & addrKnown_7; // @[LoadQueue.scala 152:41:@12881.4]
  assign _T_15022 = addrQ_7 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12882.4]
  assign conflict_7_5 = _T_15021 & _T_15022; // @[LoadQueue.scala 152:68:@12883.4]
  assign _T_15024 = entriesToCheck_7_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12885.4]
  assign _T_15025 = _T_15024 & addrKnown_7; // @[LoadQueue.scala 152:41:@12886.4]
  assign _T_15026 = addrQ_7 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12887.4]
  assign conflict_7_6 = _T_15025 & _T_15026; // @[LoadQueue.scala 152:68:@12888.4]
  assign _T_15028 = entriesToCheck_7_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12890.4]
  assign _T_15029 = _T_15028 & addrKnown_7; // @[LoadQueue.scala 152:41:@12891.4]
  assign _T_15030 = addrQ_7 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12892.4]
  assign conflict_7_7 = _T_15029 & _T_15030; // @[LoadQueue.scala 152:68:@12893.4]
  assign _T_15032 = entriesToCheck_7_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12895.4]
  assign _T_15033 = _T_15032 & addrKnown_7; // @[LoadQueue.scala 152:41:@12896.4]
  assign _T_15034 = addrQ_7 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12897.4]
  assign conflict_7_8 = _T_15033 & _T_15034; // @[LoadQueue.scala 152:68:@12898.4]
  assign _T_15036 = entriesToCheck_7_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12900.4]
  assign _T_15037 = _T_15036 & addrKnown_7; // @[LoadQueue.scala 152:41:@12901.4]
  assign _T_15038 = addrQ_7 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12902.4]
  assign conflict_7_9 = _T_15037 & _T_15038; // @[LoadQueue.scala 152:68:@12903.4]
  assign _T_15040 = entriesToCheck_7_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12905.4]
  assign _T_15041 = _T_15040 & addrKnown_7; // @[LoadQueue.scala 152:41:@12906.4]
  assign _T_15042 = addrQ_7 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12907.4]
  assign conflict_7_10 = _T_15041 & _T_15042; // @[LoadQueue.scala 152:68:@12908.4]
  assign _T_15044 = entriesToCheck_7_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12910.4]
  assign _T_15045 = _T_15044 & addrKnown_7; // @[LoadQueue.scala 152:41:@12911.4]
  assign _T_15046 = addrQ_7 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12912.4]
  assign conflict_7_11 = _T_15045 & _T_15046; // @[LoadQueue.scala 152:68:@12913.4]
  assign _T_15048 = entriesToCheck_7_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12915.4]
  assign _T_15049 = _T_15048 & addrKnown_7; // @[LoadQueue.scala 152:41:@12916.4]
  assign _T_15050 = addrQ_7 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12917.4]
  assign conflict_7_12 = _T_15049 & _T_15050; // @[LoadQueue.scala 152:68:@12918.4]
  assign _T_15052 = entriesToCheck_7_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@12920.4]
  assign _T_15053 = _T_15052 & addrKnown_7; // @[LoadQueue.scala 152:41:@12921.4]
  assign _T_15054 = addrQ_7 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@12922.4]
  assign conflict_7_13 = _T_15053 & _T_15054; // @[LoadQueue.scala 152:68:@12923.4]
  assign _T_15056 = entriesToCheck_7_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@12925.4]
  assign _T_15057 = _T_15056 & addrKnown_7; // @[LoadQueue.scala 152:41:@12926.4]
  assign _T_15058 = addrQ_7 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@12927.4]
  assign conflict_7_14 = _T_15057 & _T_15058; // @[LoadQueue.scala 152:68:@12928.4]
  assign _T_15060 = entriesToCheck_7_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@12930.4]
  assign _T_15061 = _T_15060 & addrKnown_7; // @[LoadQueue.scala 152:41:@12931.4]
  assign _T_15062 = addrQ_7 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@12932.4]
  assign conflict_7_15 = _T_15061 & _T_15062; // @[LoadQueue.scala 152:68:@12933.4]
  assign _T_15064 = entriesToCheck_8_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12935.4]
  assign _T_15065 = _T_15064 & addrKnown_8; // @[LoadQueue.scala 152:41:@12936.4]
  assign _T_15066 = addrQ_8 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12937.4]
  assign conflict_8_0 = _T_15065 & _T_15066; // @[LoadQueue.scala 152:68:@12938.4]
  assign _T_15068 = entriesToCheck_8_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12940.4]
  assign _T_15069 = _T_15068 & addrKnown_8; // @[LoadQueue.scala 152:41:@12941.4]
  assign _T_15070 = addrQ_8 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12942.4]
  assign conflict_8_1 = _T_15069 & _T_15070; // @[LoadQueue.scala 152:68:@12943.4]
  assign _T_15072 = entriesToCheck_8_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12945.4]
  assign _T_15073 = _T_15072 & addrKnown_8; // @[LoadQueue.scala 152:41:@12946.4]
  assign _T_15074 = addrQ_8 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12947.4]
  assign conflict_8_2 = _T_15073 & _T_15074; // @[LoadQueue.scala 152:68:@12948.4]
  assign _T_15076 = entriesToCheck_8_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12950.4]
  assign _T_15077 = _T_15076 & addrKnown_8; // @[LoadQueue.scala 152:41:@12951.4]
  assign _T_15078 = addrQ_8 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12952.4]
  assign conflict_8_3 = _T_15077 & _T_15078; // @[LoadQueue.scala 152:68:@12953.4]
  assign _T_15080 = entriesToCheck_8_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12955.4]
  assign _T_15081 = _T_15080 & addrKnown_8; // @[LoadQueue.scala 152:41:@12956.4]
  assign _T_15082 = addrQ_8 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12957.4]
  assign conflict_8_4 = _T_15081 & _T_15082; // @[LoadQueue.scala 152:68:@12958.4]
  assign _T_15084 = entriesToCheck_8_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12960.4]
  assign _T_15085 = _T_15084 & addrKnown_8; // @[LoadQueue.scala 152:41:@12961.4]
  assign _T_15086 = addrQ_8 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12962.4]
  assign conflict_8_5 = _T_15085 & _T_15086; // @[LoadQueue.scala 152:68:@12963.4]
  assign _T_15088 = entriesToCheck_8_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12965.4]
  assign _T_15089 = _T_15088 & addrKnown_8; // @[LoadQueue.scala 152:41:@12966.4]
  assign _T_15090 = addrQ_8 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12967.4]
  assign conflict_8_6 = _T_15089 & _T_15090; // @[LoadQueue.scala 152:68:@12968.4]
  assign _T_15092 = entriesToCheck_8_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12970.4]
  assign _T_15093 = _T_15092 & addrKnown_8; // @[LoadQueue.scala 152:41:@12971.4]
  assign _T_15094 = addrQ_8 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12972.4]
  assign conflict_8_7 = _T_15093 & _T_15094; // @[LoadQueue.scala 152:68:@12973.4]
  assign _T_15096 = entriesToCheck_8_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12975.4]
  assign _T_15097 = _T_15096 & addrKnown_8; // @[LoadQueue.scala 152:41:@12976.4]
  assign _T_15098 = addrQ_8 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12977.4]
  assign conflict_8_8 = _T_15097 & _T_15098; // @[LoadQueue.scala 152:68:@12978.4]
  assign _T_15100 = entriesToCheck_8_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12980.4]
  assign _T_15101 = _T_15100 & addrKnown_8; // @[LoadQueue.scala 152:41:@12981.4]
  assign _T_15102 = addrQ_8 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12982.4]
  assign conflict_8_9 = _T_15101 & _T_15102; // @[LoadQueue.scala 152:68:@12983.4]
  assign _T_15104 = entriesToCheck_8_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12985.4]
  assign _T_15105 = _T_15104 & addrKnown_8; // @[LoadQueue.scala 152:41:@12986.4]
  assign _T_15106 = addrQ_8 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12987.4]
  assign conflict_8_10 = _T_15105 & _T_15106; // @[LoadQueue.scala 152:68:@12988.4]
  assign _T_15108 = entriesToCheck_8_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12990.4]
  assign _T_15109 = _T_15108 & addrKnown_8; // @[LoadQueue.scala 152:41:@12991.4]
  assign _T_15110 = addrQ_8 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12992.4]
  assign conflict_8_11 = _T_15109 & _T_15110; // @[LoadQueue.scala 152:68:@12993.4]
  assign _T_15112 = entriesToCheck_8_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12995.4]
  assign _T_15113 = _T_15112 & addrKnown_8; // @[LoadQueue.scala 152:41:@12996.4]
  assign _T_15114 = addrQ_8 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12997.4]
  assign conflict_8_12 = _T_15113 & _T_15114; // @[LoadQueue.scala 152:68:@12998.4]
  assign _T_15116 = entriesToCheck_8_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@13000.4]
  assign _T_15117 = _T_15116 & addrKnown_8; // @[LoadQueue.scala 152:41:@13001.4]
  assign _T_15118 = addrQ_8 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@13002.4]
  assign conflict_8_13 = _T_15117 & _T_15118; // @[LoadQueue.scala 152:68:@13003.4]
  assign _T_15120 = entriesToCheck_8_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@13005.4]
  assign _T_15121 = _T_15120 & addrKnown_8; // @[LoadQueue.scala 152:41:@13006.4]
  assign _T_15122 = addrQ_8 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@13007.4]
  assign conflict_8_14 = _T_15121 & _T_15122; // @[LoadQueue.scala 152:68:@13008.4]
  assign _T_15124 = entriesToCheck_8_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@13010.4]
  assign _T_15125 = _T_15124 & addrKnown_8; // @[LoadQueue.scala 152:41:@13011.4]
  assign _T_15126 = addrQ_8 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@13012.4]
  assign conflict_8_15 = _T_15125 & _T_15126; // @[LoadQueue.scala 152:68:@13013.4]
  assign _T_15128 = entriesToCheck_9_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@13015.4]
  assign _T_15129 = _T_15128 & addrKnown_9; // @[LoadQueue.scala 152:41:@13016.4]
  assign _T_15130 = addrQ_9 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@13017.4]
  assign conflict_9_0 = _T_15129 & _T_15130; // @[LoadQueue.scala 152:68:@13018.4]
  assign _T_15132 = entriesToCheck_9_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@13020.4]
  assign _T_15133 = _T_15132 & addrKnown_9; // @[LoadQueue.scala 152:41:@13021.4]
  assign _T_15134 = addrQ_9 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@13022.4]
  assign conflict_9_1 = _T_15133 & _T_15134; // @[LoadQueue.scala 152:68:@13023.4]
  assign _T_15136 = entriesToCheck_9_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@13025.4]
  assign _T_15137 = _T_15136 & addrKnown_9; // @[LoadQueue.scala 152:41:@13026.4]
  assign _T_15138 = addrQ_9 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@13027.4]
  assign conflict_9_2 = _T_15137 & _T_15138; // @[LoadQueue.scala 152:68:@13028.4]
  assign _T_15140 = entriesToCheck_9_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@13030.4]
  assign _T_15141 = _T_15140 & addrKnown_9; // @[LoadQueue.scala 152:41:@13031.4]
  assign _T_15142 = addrQ_9 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@13032.4]
  assign conflict_9_3 = _T_15141 & _T_15142; // @[LoadQueue.scala 152:68:@13033.4]
  assign _T_15144 = entriesToCheck_9_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@13035.4]
  assign _T_15145 = _T_15144 & addrKnown_9; // @[LoadQueue.scala 152:41:@13036.4]
  assign _T_15146 = addrQ_9 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@13037.4]
  assign conflict_9_4 = _T_15145 & _T_15146; // @[LoadQueue.scala 152:68:@13038.4]
  assign _T_15148 = entriesToCheck_9_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@13040.4]
  assign _T_15149 = _T_15148 & addrKnown_9; // @[LoadQueue.scala 152:41:@13041.4]
  assign _T_15150 = addrQ_9 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@13042.4]
  assign conflict_9_5 = _T_15149 & _T_15150; // @[LoadQueue.scala 152:68:@13043.4]
  assign _T_15152 = entriesToCheck_9_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@13045.4]
  assign _T_15153 = _T_15152 & addrKnown_9; // @[LoadQueue.scala 152:41:@13046.4]
  assign _T_15154 = addrQ_9 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@13047.4]
  assign conflict_9_6 = _T_15153 & _T_15154; // @[LoadQueue.scala 152:68:@13048.4]
  assign _T_15156 = entriesToCheck_9_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@13050.4]
  assign _T_15157 = _T_15156 & addrKnown_9; // @[LoadQueue.scala 152:41:@13051.4]
  assign _T_15158 = addrQ_9 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@13052.4]
  assign conflict_9_7 = _T_15157 & _T_15158; // @[LoadQueue.scala 152:68:@13053.4]
  assign _T_15160 = entriesToCheck_9_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@13055.4]
  assign _T_15161 = _T_15160 & addrKnown_9; // @[LoadQueue.scala 152:41:@13056.4]
  assign _T_15162 = addrQ_9 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@13057.4]
  assign conflict_9_8 = _T_15161 & _T_15162; // @[LoadQueue.scala 152:68:@13058.4]
  assign _T_15164 = entriesToCheck_9_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@13060.4]
  assign _T_15165 = _T_15164 & addrKnown_9; // @[LoadQueue.scala 152:41:@13061.4]
  assign _T_15166 = addrQ_9 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@13062.4]
  assign conflict_9_9 = _T_15165 & _T_15166; // @[LoadQueue.scala 152:68:@13063.4]
  assign _T_15168 = entriesToCheck_9_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@13065.4]
  assign _T_15169 = _T_15168 & addrKnown_9; // @[LoadQueue.scala 152:41:@13066.4]
  assign _T_15170 = addrQ_9 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@13067.4]
  assign conflict_9_10 = _T_15169 & _T_15170; // @[LoadQueue.scala 152:68:@13068.4]
  assign _T_15172 = entriesToCheck_9_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@13070.4]
  assign _T_15173 = _T_15172 & addrKnown_9; // @[LoadQueue.scala 152:41:@13071.4]
  assign _T_15174 = addrQ_9 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@13072.4]
  assign conflict_9_11 = _T_15173 & _T_15174; // @[LoadQueue.scala 152:68:@13073.4]
  assign _T_15176 = entriesToCheck_9_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@13075.4]
  assign _T_15177 = _T_15176 & addrKnown_9; // @[LoadQueue.scala 152:41:@13076.4]
  assign _T_15178 = addrQ_9 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@13077.4]
  assign conflict_9_12 = _T_15177 & _T_15178; // @[LoadQueue.scala 152:68:@13078.4]
  assign _T_15180 = entriesToCheck_9_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@13080.4]
  assign _T_15181 = _T_15180 & addrKnown_9; // @[LoadQueue.scala 152:41:@13081.4]
  assign _T_15182 = addrQ_9 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@13082.4]
  assign conflict_9_13 = _T_15181 & _T_15182; // @[LoadQueue.scala 152:68:@13083.4]
  assign _T_15184 = entriesToCheck_9_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@13085.4]
  assign _T_15185 = _T_15184 & addrKnown_9; // @[LoadQueue.scala 152:41:@13086.4]
  assign _T_15186 = addrQ_9 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@13087.4]
  assign conflict_9_14 = _T_15185 & _T_15186; // @[LoadQueue.scala 152:68:@13088.4]
  assign _T_15188 = entriesToCheck_9_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@13090.4]
  assign _T_15189 = _T_15188 & addrKnown_9; // @[LoadQueue.scala 152:41:@13091.4]
  assign _T_15190 = addrQ_9 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@13092.4]
  assign conflict_9_15 = _T_15189 & _T_15190; // @[LoadQueue.scala 152:68:@13093.4]
  assign _T_15192 = entriesToCheck_10_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@13095.4]
  assign _T_15193 = _T_15192 & addrKnown_10; // @[LoadQueue.scala 152:41:@13096.4]
  assign _T_15194 = addrQ_10 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@13097.4]
  assign conflict_10_0 = _T_15193 & _T_15194; // @[LoadQueue.scala 152:68:@13098.4]
  assign _T_15196 = entriesToCheck_10_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@13100.4]
  assign _T_15197 = _T_15196 & addrKnown_10; // @[LoadQueue.scala 152:41:@13101.4]
  assign _T_15198 = addrQ_10 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@13102.4]
  assign conflict_10_1 = _T_15197 & _T_15198; // @[LoadQueue.scala 152:68:@13103.4]
  assign _T_15200 = entriesToCheck_10_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@13105.4]
  assign _T_15201 = _T_15200 & addrKnown_10; // @[LoadQueue.scala 152:41:@13106.4]
  assign _T_15202 = addrQ_10 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@13107.4]
  assign conflict_10_2 = _T_15201 & _T_15202; // @[LoadQueue.scala 152:68:@13108.4]
  assign _T_15204 = entriesToCheck_10_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@13110.4]
  assign _T_15205 = _T_15204 & addrKnown_10; // @[LoadQueue.scala 152:41:@13111.4]
  assign _T_15206 = addrQ_10 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@13112.4]
  assign conflict_10_3 = _T_15205 & _T_15206; // @[LoadQueue.scala 152:68:@13113.4]
  assign _T_15208 = entriesToCheck_10_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@13115.4]
  assign _T_15209 = _T_15208 & addrKnown_10; // @[LoadQueue.scala 152:41:@13116.4]
  assign _T_15210 = addrQ_10 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@13117.4]
  assign conflict_10_4 = _T_15209 & _T_15210; // @[LoadQueue.scala 152:68:@13118.4]
  assign _T_15212 = entriesToCheck_10_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@13120.4]
  assign _T_15213 = _T_15212 & addrKnown_10; // @[LoadQueue.scala 152:41:@13121.4]
  assign _T_15214 = addrQ_10 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@13122.4]
  assign conflict_10_5 = _T_15213 & _T_15214; // @[LoadQueue.scala 152:68:@13123.4]
  assign _T_15216 = entriesToCheck_10_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@13125.4]
  assign _T_15217 = _T_15216 & addrKnown_10; // @[LoadQueue.scala 152:41:@13126.4]
  assign _T_15218 = addrQ_10 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@13127.4]
  assign conflict_10_6 = _T_15217 & _T_15218; // @[LoadQueue.scala 152:68:@13128.4]
  assign _T_15220 = entriesToCheck_10_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@13130.4]
  assign _T_15221 = _T_15220 & addrKnown_10; // @[LoadQueue.scala 152:41:@13131.4]
  assign _T_15222 = addrQ_10 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@13132.4]
  assign conflict_10_7 = _T_15221 & _T_15222; // @[LoadQueue.scala 152:68:@13133.4]
  assign _T_15224 = entriesToCheck_10_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@13135.4]
  assign _T_15225 = _T_15224 & addrKnown_10; // @[LoadQueue.scala 152:41:@13136.4]
  assign _T_15226 = addrQ_10 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@13137.4]
  assign conflict_10_8 = _T_15225 & _T_15226; // @[LoadQueue.scala 152:68:@13138.4]
  assign _T_15228 = entriesToCheck_10_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@13140.4]
  assign _T_15229 = _T_15228 & addrKnown_10; // @[LoadQueue.scala 152:41:@13141.4]
  assign _T_15230 = addrQ_10 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@13142.4]
  assign conflict_10_9 = _T_15229 & _T_15230; // @[LoadQueue.scala 152:68:@13143.4]
  assign _T_15232 = entriesToCheck_10_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@13145.4]
  assign _T_15233 = _T_15232 & addrKnown_10; // @[LoadQueue.scala 152:41:@13146.4]
  assign _T_15234 = addrQ_10 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@13147.4]
  assign conflict_10_10 = _T_15233 & _T_15234; // @[LoadQueue.scala 152:68:@13148.4]
  assign _T_15236 = entriesToCheck_10_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@13150.4]
  assign _T_15237 = _T_15236 & addrKnown_10; // @[LoadQueue.scala 152:41:@13151.4]
  assign _T_15238 = addrQ_10 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@13152.4]
  assign conflict_10_11 = _T_15237 & _T_15238; // @[LoadQueue.scala 152:68:@13153.4]
  assign _T_15240 = entriesToCheck_10_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@13155.4]
  assign _T_15241 = _T_15240 & addrKnown_10; // @[LoadQueue.scala 152:41:@13156.4]
  assign _T_15242 = addrQ_10 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@13157.4]
  assign conflict_10_12 = _T_15241 & _T_15242; // @[LoadQueue.scala 152:68:@13158.4]
  assign _T_15244 = entriesToCheck_10_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@13160.4]
  assign _T_15245 = _T_15244 & addrKnown_10; // @[LoadQueue.scala 152:41:@13161.4]
  assign _T_15246 = addrQ_10 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@13162.4]
  assign conflict_10_13 = _T_15245 & _T_15246; // @[LoadQueue.scala 152:68:@13163.4]
  assign _T_15248 = entriesToCheck_10_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@13165.4]
  assign _T_15249 = _T_15248 & addrKnown_10; // @[LoadQueue.scala 152:41:@13166.4]
  assign _T_15250 = addrQ_10 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@13167.4]
  assign conflict_10_14 = _T_15249 & _T_15250; // @[LoadQueue.scala 152:68:@13168.4]
  assign _T_15252 = entriesToCheck_10_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@13170.4]
  assign _T_15253 = _T_15252 & addrKnown_10; // @[LoadQueue.scala 152:41:@13171.4]
  assign _T_15254 = addrQ_10 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@13172.4]
  assign conflict_10_15 = _T_15253 & _T_15254; // @[LoadQueue.scala 152:68:@13173.4]
  assign _T_15256 = entriesToCheck_11_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@13175.4]
  assign _T_15257 = _T_15256 & addrKnown_11; // @[LoadQueue.scala 152:41:@13176.4]
  assign _T_15258 = addrQ_11 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@13177.4]
  assign conflict_11_0 = _T_15257 & _T_15258; // @[LoadQueue.scala 152:68:@13178.4]
  assign _T_15260 = entriesToCheck_11_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@13180.4]
  assign _T_15261 = _T_15260 & addrKnown_11; // @[LoadQueue.scala 152:41:@13181.4]
  assign _T_15262 = addrQ_11 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@13182.4]
  assign conflict_11_1 = _T_15261 & _T_15262; // @[LoadQueue.scala 152:68:@13183.4]
  assign _T_15264 = entriesToCheck_11_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@13185.4]
  assign _T_15265 = _T_15264 & addrKnown_11; // @[LoadQueue.scala 152:41:@13186.4]
  assign _T_15266 = addrQ_11 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@13187.4]
  assign conflict_11_2 = _T_15265 & _T_15266; // @[LoadQueue.scala 152:68:@13188.4]
  assign _T_15268 = entriesToCheck_11_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@13190.4]
  assign _T_15269 = _T_15268 & addrKnown_11; // @[LoadQueue.scala 152:41:@13191.4]
  assign _T_15270 = addrQ_11 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@13192.4]
  assign conflict_11_3 = _T_15269 & _T_15270; // @[LoadQueue.scala 152:68:@13193.4]
  assign _T_15272 = entriesToCheck_11_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@13195.4]
  assign _T_15273 = _T_15272 & addrKnown_11; // @[LoadQueue.scala 152:41:@13196.4]
  assign _T_15274 = addrQ_11 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@13197.4]
  assign conflict_11_4 = _T_15273 & _T_15274; // @[LoadQueue.scala 152:68:@13198.4]
  assign _T_15276 = entriesToCheck_11_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@13200.4]
  assign _T_15277 = _T_15276 & addrKnown_11; // @[LoadQueue.scala 152:41:@13201.4]
  assign _T_15278 = addrQ_11 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@13202.4]
  assign conflict_11_5 = _T_15277 & _T_15278; // @[LoadQueue.scala 152:68:@13203.4]
  assign _T_15280 = entriesToCheck_11_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@13205.4]
  assign _T_15281 = _T_15280 & addrKnown_11; // @[LoadQueue.scala 152:41:@13206.4]
  assign _T_15282 = addrQ_11 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@13207.4]
  assign conflict_11_6 = _T_15281 & _T_15282; // @[LoadQueue.scala 152:68:@13208.4]
  assign _T_15284 = entriesToCheck_11_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@13210.4]
  assign _T_15285 = _T_15284 & addrKnown_11; // @[LoadQueue.scala 152:41:@13211.4]
  assign _T_15286 = addrQ_11 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@13212.4]
  assign conflict_11_7 = _T_15285 & _T_15286; // @[LoadQueue.scala 152:68:@13213.4]
  assign _T_15288 = entriesToCheck_11_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@13215.4]
  assign _T_15289 = _T_15288 & addrKnown_11; // @[LoadQueue.scala 152:41:@13216.4]
  assign _T_15290 = addrQ_11 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@13217.4]
  assign conflict_11_8 = _T_15289 & _T_15290; // @[LoadQueue.scala 152:68:@13218.4]
  assign _T_15292 = entriesToCheck_11_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@13220.4]
  assign _T_15293 = _T_15292 & addrKnown_11; // @[LoadQueue.scala 152:41:@13221.4]
  assign _T_15294 = addrQ_11 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@13222.4]
  assign conflict_11_9 = _T_15293 & _T_15294; // @[LoadQueue.scala 152:68:@13223.4]
  assign _T_15296 = entriesToCheck_11_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@13225.4]
  assign _T_15297 = _T_15296 & addrKnown_11; // @[LoadQueue.scala 152:41:@13226.4]
  assign _T_15298 = addrQ_11 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@13227.4]
  assign conflict_11_10 = _T_15297 & _T_15298; // @[LoadQueue.scala 152:68:@13228.4]
  assign _T_15300 = entriesToCheck_11_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@13230.4]
  assign _T_15301 = _T_15300 & addrKnown_11; // @[LoadQueue.scala 152:41:@13231.4]
  assign _T_15302 = addrQ_11 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@13232.4]
  assign conflict_11_11 = _T_15301 & _T_15302; // @[LoadQueue.scala 152:68:@13233.4]
  assign _T_15304 = entriesToCheck_11_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@13235.4]
  assign _T_15305 = _T_15304 & addrKnown_11; // @[LoadQueue.scala 152:41:@13236.4]
  assign _T_15306 = addrQ_11 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@13237.4]
  assign conflict_11_12 = _T_15305 & _T_15306; // @[LoadQueue.scala 152:68:@13238.4]
  assign _T_15308 = entriesToCheck_11_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@13240.4]
  assign _T_15309 = _T_15308 & addrKnown_11; // @[LoadQueue.scala 152:41:@13241.4]
  assign _T_15310 = addrQ_11 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@13242.4]
  assign conflict_11_13 = _T_15309 & _T_15310; // @[LoadQueue.scala 152:68:@13243.4]
  assign _T_15312 = entriesToCheck_11_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@13245.4]
  assign _T_15313 = _T_15312 & addrKnown_11; // @[LoadQueue.scala 152:41:@13246.4]
  assign _T_15314 = addrQ_11 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@13247.4]
  assign conflict_11_14 = _T_15313 & _T_15314; // @[LoadQueue.scala 152:68:@13248.4]
  assign _T_15316 = entriesToCheck_11_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@13250.4]
  assign _T_15317 = _T_15316 & addrKnown_11; // @[LoadQueue.scala 152:41:@13251.4]
  assign _T_15318 = addrQ_11 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@13252.4]
  assign conflict_11_15 = _T_15317 & _T_15318; // @[LoadQueue.scala 152:68:@13253.4]
  assign _T_15320 = entriesToCheck_12_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@13255.4]
  assign _T_15321 = _T_15320 & addrKnown_12; // @[LoadQueue.scala 152:41:@13256.4]
  assign _T_15322 = addrQ_12 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@13257.4]
  assign conflict_12_0 = _T_15321 & _T_15322; // @[LoadQueue.scala 152:68:@13258.4]
  assign _T_15324 = entriesToCheck_12_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@13260.4]
  assign _T_15325 = _T_15324 & addrKnown_12; // @[LoadQueue.scala 152:41:@13261.4]
  assign _T_15326 = addrQ_12 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@13262.4]
  assign conflict_12_1 = _T_15325 & _T_15326; // @[LoadQueue.scala 152:68:@13263.4]
  assign _T_15328 = entriesToCheck_12_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@13265.4]
  assign _T_15329 = _T_15328 & addrKnown_12; // @[LoadQueue.scala 152:41:@13266.4]
  assign _T_15330 = addrQ_12 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@13267.4]
  assign conflict_12_2 = _T_15329 & _T_15330; // @[LoadQueue.scala 152:68:@13268.4]
  assign _T_15332 = entriesToCheck_12_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@13270.4]
  assign _T_15333 = _T_15332 & addrKnown_12; // @[LoadQueue.scala 152:41:@13271.4]
  assign _T_15334 = addrQ_12 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@13272.4]
  assign conflict_12_3 = _T_15333 & _T_15334; // @[LoadQueue.scala 152:68:@13273.4]
  assign _T_15336 = entriesToCheck_12_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@13275.4]
  assign _T_15337 = _T_15336 & addrKnown_12; // @[LoadQueue.scala 152:41:@13276.4]
  assign _T_15338 = addrQ_12 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@13277.4]
  assign conflict_12_4 = _T_15337 & _T_15338; // @[LoadQueue.scala 152:68:@13278.4]
  assign _T_15340 = entriesToCheck_12_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@13280.4]
  assign _T_15341 = _T_15340 & addrKnown_12; // @[LoadQueue.scala 152:41:@13281.4]
  assign _T_15342 = addrQ_12 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@13282.4]
  assign conflict_12_5 = _T_15341 & _T_15342; // @[LoadQueue.scala 152:68:@13283.4]
  assign _T_15344 = entriesToCheck_12_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@13285.4]
  assign _T_15345 = _T_15344 & addrKnown_12; // @[LoadQueue.scala 152:41:@13286.4]
  assign _T_15346 = addrQ_12 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@13287.4]
  assign conflict_12_6 = _T_15345 & _T_15346; // @[LoadQueue.scala 152:68:@13288.4]
  assign _T_15348 = entriesToCheck_12_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@13290.4]
  assign _T_15349 = _T_15348 & addrKnown_12; // @[LoadQueue.scala 152:41:@13291.4]
  assign _T_15350 = addrQ_12 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@13292.4]
  assign conflict_12_7 = _T_15349 & _T_15350; // @[LoadQueue.scala 152:68:@13293.4]
  assign _T_15352 = entriesToCheck_12_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@13295.4]
  assign _T_15353 = _T_15352 & addrKnown_12; // @[LoadQueue.scala 152:41:@13296.4]
  assign _T_15354 = addrQ_12 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@13297.4]
  assign conflict_12_8 = _T_15353 & _T_15354; // @[LoadQueue.scala 152:68:@13298.4]
  assign _T_15356 = entriesToCheck_12_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@13300.4]
  assign _T_15357 = _T_15356 & addrKnown_12; // @[LoadQueue.scala 152:41:@13301.4]
  assign _T_15358 = addrQ_12 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@13302.4]
  assign conflict_12_9 = _T_15357 & _T_15358; // @[LoadQueue.scala 152:68:@13303.4]
  assign _T_15360 = entriesToCheck_12_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@13305.4]
  assign _T_15361 = _T_15360 & addrKnown_12; // @[LoadQueue.scala 152:41:@13306.4]
  assign _T_15362 = addrQ_12 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@13307.4]
  assign conflict_12_10 = _T_15361 & _T_15362; // @[LoadQueue.scala 152:68:@13308.4]
  assign _T_15364 = entriesToCheck_12_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@13310.4]
  assign _T_15365 = _T_15364 & addrKnown_12; // @[LoadQueue.scala 152:41:@13311.4]
  assign _T_15366 = addrQ_12 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@13312.4]
  assign conflict_12_11 = _T_15365 & _T_15366; // @[LoadQueue.scala 152:68:@13313.4]
  assign _T_15368 = entriesToCheck_12_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@13315.4]
  assign _T_15369 = _T_15368 & addrKnown_12; // @[LoadQueue.scala 152:41:@13316.4]
  assign _T_15370 = addrQ_12 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@13317.4]
  assign conflict_12_12 = _T_15369 & _T_15370; // @[LoadQueue.scala 152:68:@13318.4]
  assign _T_15372 = entriesToCheck_12_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@13320.4]
  assign _T_15373 = _T_15372 & addrKnown_12; // @[LoadQueue.scala 152:41:@13321.4]
  assign _T_15374 = addrQ_12 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@13322.4]
  assign conflict_12_13 = _T_15373 & _T_15374; // @[LoadQueue.scala 152:68:@13323.4]
  assign _T_15376 = entriesToCheck_12_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@13325.4]
  assign _T_15377 = _T_15376 & addrKnown_12; // @[LoadQueue.scala 152:41:@13326.4]
  assign _T_15378 = addrQ_12 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@13327.4]
  assign conflict_12_14 = _T_15377 & _T_15378; // @[LoadQueue.scala 152:68:@13328.4]
  assign _T_15380 = entriesToCheck_12_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@13330.4]
  assign _T_15381 = _T_15380 & addrKnown_12; // @[LoadQueue.scala 152:41:@13331.4]
  assign _T_15382 = addrQ_12 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@13332.4]
  assign conflict_12_15 = _T_15381 & _T_15382; // @[LoadQueue.scala 152:68:@13333.4]
  assign _T_15384 = entriesToCheck_13_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@13335.4]
  assign _T_15385 = _T_15384 & addrKnown_13; // @[LoadQueue.scala 152:41:@13336.4]
  assign _T_15386 = addrQ_13 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@13337.4]
  assign conflict_13_0 = _T_15385 & _T_15386; // @[LoadQueue.scala 152:68:@13338.4]
  assign _T_15388 = entriesToCheck_13_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@13340.4]
  assign _T_15389 = _T_15388 & addrKnown_13; // @[LoadQueue.scala 152:41:@13341.4]
  assign _T_15390 = addrQ_13 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@13342.4]
  assign conflict_13_1 = _T_15389 & _T_15390; // @[LoadQueue.scala 152:68:@13343.4]
  assign _T_15392 = entriesToCheck_13_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@13345.4]
  assign _T_15393 = _T_15392 & addrKnown_13; // @[LoadQueue.scala 152:41:@13346.4]
  assign _T_15394 = addrQ_13 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@13347.4]
  assign conflict_13_2 = _T_15393 & _T_15394; // @[LoadQueue.scala 152:68:@13348.4]
  assign _T_15396 = entriesToCheck_13_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@13350.4]
  assign _T_15397 = _T_15396 & addrKnown_13; // @[LoadQueue.scala 152:41:@13351.4]
  assign _T_15398 = addrQ_13 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@13352.4]
  assign conflict_13_3 = _T_15397 & _T_15398; // @[LoadQueue.scala 152:68:@13353.4]
  assign _T_15400 = entriesToCheck_13_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@13355.4]
  assign _T_15401 = _T_15400 & addrKnown_13; // @[LoadQueue.scala 152:41:@13356.4]
  assign _T_15402 = addrQ_13 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@13357.4]
  assign conflict_13_4 = _T_15401 & _T_15402; // @[LoadQueue.scala 152:68:@13358.4]
  assign _T_15404 = entriesToCheck_13_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@13360.4]
  assign _T_15405 = _T_15404 & addrKnown_13; // @[LoadQueue.scala 152:41:@13361.4]
  assign _T_15406 = addrQ_13 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@13362.4]
  assign conflict_13_5 = _T_15405 & _T_15406; // @[LoadQueue.scala 152:68:@13363.4]
  assign _T_15408 = entriesToCheck_13_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@13365.4]
  assign _T_15409 = _T_15408 & addrKnown_13; // @[LoadQueue.scala 152:41:@13366.4]
  assign _T_15410 = addrQ_13 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@13367.4]
  assign conflict_13_6 = _T_15409 & _T_15410; // @[LoadQueue.scala 152:68:@13368.4]
  assign _T_15412 = entriesToCheck_13_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@13370.4]
  assign _T_15413 = _T_15412 & addrKnown_13; // @[LoadQueue.scala 152:41:@13371.4]
  assign _T_15414 = addrQ_13 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@13372.4]
  assign conflict_13_7 = _T_15413 & _T_15414; // @[LoadQueue.scala 152:68:@13373.4]
  assign _T_15416 = entriesToCheck_13_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@13375.4]
  assign _T_15417 = _T_15416 & addrKnown_13; // @[LoadQueue.scala 152:41:@13376.4]
  assign _T_15418 = addrQ_13 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@13377.4]
  assign conflict_13_8 = _T_15417 & _T_15418; // @[LoadQueue.scala 152:68:@13378.4]
  assign _T_15420 = entriesToCheck_13_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@13380.4]
  assign _T_15421 = _T_15420 & addrKnown_13; // @[LoadQueue.scala 152:41:@13381.4]
  assign _T_15422 = addrQ_13 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@13382.4]
  assign conflict_13_9 = _T_15421 & _T_15422; // @[LoadQueue.scala 152:68:@13383.4]
  assign _T_15424 = entriesToCheck_13_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@13385.4]
  assign _T_15425 = _T_15424 & addrKnown_13; // @[LoadQueue.scala 152:41:@13386.4]
  assign _T_15426 = addrQ_13 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@13387.4]
  assign conflict_13_10 = _T_15425 & _T_15426; // @[LoadQueue.scala 152:68:@13388.4]
  assign _T_15428 = entriesToCheck_13_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@13390.4]
  assign _T_15429 = _T_15428 & addrKnown_13; // @[LoadQueue.scala 152:41:@13391.4]
  assign _T_15430 = addrQ_13 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@13392.4]
  assign conflict_13_11 = _T_15429 & _T_15430; // @[LoadQueue.scala 152:68:@13393.4]
  assign _T_15432 = entriesToCheck_13_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@13395.4]
  assign _T_15433 = _T_15432 & addrKnown_13; // @[LoadQueue.scala 152:41:@13396.4]
  assign _T_15434 = addrQ_13 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@13397.4]
  assign conflict_13_12 = _T_15433 & _T_15434; // @[LoadQueue.scala 152:68:@13398.4]
  assign _T_15436 = entriesToCheck_13_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@13400.4]
  assign _T_15437 = _T_15436 & addrKnown_13; // @[LoadQueue.scala 152:41:@13401.4]
  assign _T_15438 = addrQ_13 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@13402.4]
  assign conflict_13_13 = _T_15437 & _T_15438; // @[LoadQueue.scala 152:68:@13403.4]
  assign _T_15440 = entriesToCheck_13_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@13405.4]
  assign _T_15441 = _T_15440 & addrKnown_13; // @[LoadQueue.scala 152:41:@13406.4]
  assign _T_15442 = addrQ_13 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@13407.4]
  assign conflict_13_14 = _T_15441 & _T_15442; // @[LoadQueue.scala 152:68:@13408.4]
  assign _T_15444 = entriesToCheck_13_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@13410.4]
  assign _T_15445 = _T_15444 & addrKnown_13; // @[LoadQueue.scala 152:41:@13411.4]
  assign _T_15446 = addrQ_13 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@13412.4]
  assign conflict_13_15 = _T_15445 & _T_15446; // @[LoadQueue.scala 152:68:@13413.4]
  assign _T_15448 = entriesToCheck_14_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@13415.4]
  assign _T_15449 = _T_15448 & addrKnown_14; // @[LoadQueue.scala 152:41:@13416.4]
  assign _T_15450 = addrQ_14 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@13417.4]
  assign conflict_14_0 = _T_15449 & _T_15450; // @[LoadQueue.scala 152:68:@13418.4]
  assign _T_15452 = entriesToCheck_14_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@13420.4]
  assign _T_15453 = _T_15452 & addrKnown_14; // @[LoadQueue.scala 152:41:@13421.4]
  assign _T_15454 = addrQ_14 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@13422.4]
  assign conflict_14_1 = _T_15453 & _T_15454; // @[LoadQueue.scala 152:68:@13423.4]
  assign _T_15456 = entriesToCheck_14_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@13425.4]
  assign _T_15457 = _T_15456 & addrKnown_14; // @[LoadQueue.scala 152:41:@13426.4]
  assign _T_15458 = addrQ_14 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@13427.4]
  assign conflict_14_2 = _T_15457 & _T_15458; // @[LoadQueue.scala 152:68:@13428.4]
  assign _T_15460 = entriesToCheck_14_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@13430.4]
  assign _T_15461 = _T_15460 & addrKnown_14; // @[LoadQueue.scala 152:41:@13431.4]
  assign _T_15462 = addrQ_14 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@13432.4]
  assign conflict_14_3 = _T_15461 & _T_15462; // @[LoadQueue.scala 152:68:@13433.4]
  assign _T_15464 = entriesToCheck_14_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@13435.4]
  assign _T_15465 = _T_15464 & addrKnown_14; // @[LoadQueue.scala 152:41:@13436.4]
  assign _T_15466 = addrQ_14 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@13437.4]
  assign conflict_14_4 = _T_15465 & _T_15466; // @[LoadQueue.scala 152:68:@13438.4]
  assign _T_15468 = entriesToCheck_14_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@13440.4]
  assign _T_15469 = _T_15468 & addrKnown_14; // @[LoadQueue.scala 152:41:@13441.4]
  assign _T_15470 = addrQ_14 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@13442.4]
  assign conflict_14_5 = _T_15469 & _T_15470; // @[LoadQueue.scala 152:68:@13443.4]
  assign _T_15472 = entriesToCheck_14_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@13445.4]
  assign _T_15473 = _T_15472 & addrKnown_14; // @[LoadQueue.scala 152:41:@13446.4]
  assign _T_15474 = addrQ_14 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@13447.4]
  assign conflict_14_6 = _T_15473 & _T_15474; // @[LoadQueue.scala 152:68:@13448.4]
  assign _T_15476 = entriesToCheck_14_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@13450.4]
  assign _T_15477 = _T_15476 & addrKnown_14; // @[LoadQueue.scala 152:41:@13451.4]
  assign _T_15478 = addrQ_14 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@13452.4]
  assign conflict_14_7 = _T_15477 & _T_15478; // @[LoadQueue.scala 152:68:@13453.4]
  assign _T_15480 = entriesToCheck_14_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@13455.4]
  assign _T_15481 = _T_15480 & addrKnown_14; // @[LoadQueue.scala 152:41:@13456.4]
  assign _T_15482 = addrQ_14 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@13457.4]
  assign conflict_14_8 = _T_15481 & _T_15482; // @[LoadQueue.scala 152:68:@13458.4]
  assign _T_15484 = entriesToCheck_14_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@13460.4]
  assign _T_15485 = _T_15484 & addrKnown_14; // @[LoadQueue.scala 152:41:@13461.4]
  assign _T_15486 = addrQ_14 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@13462.4]
  assign conflict_14_9 = _T_15485 & _T_15486; // @[LoadQueue.scala 152:68:@13463.4]
  assign _T_15488 = entriesToCheck_14_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@13465.4]
  assign _T_15489 = _T_15488 & addrKnown_14; // @[LoadQueue.scala 152:41:@13466.4]
  assign _T_15490 = addrQ_14 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@13467.4]
  assign conflict_14_10 = _T_15489 & _T_15490; // @[LoadQueue.scala 152:68:@13468.4]
  assign _T_15492 = entriesToCheck_14_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@13470.4]
  assign _T_15493 = _T_15492 & addrKnown_14; // @[LoadQueue.scala 152:41:@13471.4]
  assign _T_15494 = addrQ_14 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@13472.4]
  assign conflict_14_11 = _T_15493 & _T_15494; // @[LoadQueue.scala 152:68:@13473.4]
  assign _T_15496 = entriesToCheck_14_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@13475.4]
  assign _T_15497 = _T_15496 & addrKnown_14; // @[LoadQueue.scala 152:41:@13476.4]
  assign _T_15498 = addrQ_14 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@13477.4]
  assign conflict_14_12 = _T_15497 & _T_15498; // @[LoadQueue.scala 152:68:@13478.4]
  assign _T_15500 = entriesToCheck_14_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@13480.4]
  assign _T_15501 = _T_15500 & addrKnown_14; // @[LoadQueue.scala 152:41:@13481.4]
  assign _T_15502 = addrQ_14 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@13482.4]
  assign conflict_14_13 = _T_15501 & _T_15502; // @[LoadQueue.scala 152:68:@13483.4]
  assign _T_15504 = entriesToCheck_14_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@13485.4]
  assign _T_15505 = _T_15504 & addrKnown_14; // @[LoadQueue.scala 152:41:@13486.4]
  assign _T_15506 = addrQ_14 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@13487.4]
  assign conflict_14_14 = _T_15505 & _T_15506; // @[LoadQueue.scala 152:68:@13488.4]
  assign _T_15508 = entriesToCheck_14_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@13490.4]
  assign _T_15509 = _T_15508 & addrKnown_14; // @[LoadQueue.scala 152:41:@13491.4]
  assign _T_15510 = addrQ_14 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@13492.4]
  assign conflict_14_15 = _T_15509 & _T_15510; // @[LoadQueue.scala 152:68:@13493.4]
  assign _T_15512 = entriesToCheck_15_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@13495.4]
  assign _T_15513 = _T_15512 & addrKnown_15; // @[LoadQueue.scala 152:41:@13496.4]
  assign _T_15514 = addrQ_15 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@13497.4]
  assign conflict_15_0 = _T_15513 & _T_15514; // @[LoadQueue.scala 152:68:@13498.4]
  assign _T_15516 = entriesToCheck_15_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@13500.4]
  assign _T_15517 = _T_15516 & addrKnown_15; // @[LoadQueue.scala 152:41:@13501.4]
  assign _T_15518 = addrQ_15 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@13502.4]
  assign conflict_15_1 = _T_15517 & _T_15518; // @[LoadQueue.scala 152:68:@13503.4]
  assign _T_15520 = entriesToCheck_15_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@13505.4]
  assign _T_15521 = _T_15520 & addrKnown_15; // @[LoadQueue.scala 152:41:@13506.4]
  assign _T_15522 = addrQ_15 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@13507.4]
  assign conflict_15_2 = _T_15521 & _T_15522; // @[LoadQueue.scala 152:68:@13508.4]
  assign _T_15524 = entriesToCheck_15_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@13510.4]
  assign _T_15525 = _T_15524 & addrKnown_15; // @[LoadQueue.scala 152:41:@13511.4]
  assign _T_15526 = addrQ_15 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@13512.4]
  assign conflict_15_3 = _T_15525 & _T_15526; // @[LoadQueue.scala 152:68:@13513.4]
  assign _T_15528 = entriesToCheck_15_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@13515.4]
  assign _T_15529 = _T_15528 & addrKnown_15; // @[LoadQueue.scala 152:41:@13516.4]
  assign _T_15530 = addrQ_15 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@13517.4]
  assign conflict_15_4 = _T_15529 & _T_15530; // @[LoadQueue.scala 152:68:@13518.4]
  assign _T_15532 = entriesToCheck_15_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@13520.4]
  assign _T_15533 = _T_15532 & addrKnown_15; // @[LoadQueue.scala 152:41:@13521.4]
  assign _T_15534 = addrQ_15 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@13522.4]
  assign conflict_15_5 = _T_15533 & _T_15534; // @[LoadQueue.scala 152:68:@13523.4]
  assign _T_15536 = entriesToCheck_15_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@13525.4]
  assign _T_15537 = _T_15536 & addrKnown_15; // @[LoadQueue.scala 152:41:@13526.4]
  assign _T_15538 = addrQ_15 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@13527.4]
  assign conflict_15_6 = _T_15537 & _T_15538; // @[LoadQueue.scala 152:68:@13528.4]
  assign _T_15540 = entriesToCheck_15_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@13530.4]
  assign _T_15541 = _T_15540 & addrKnown_15; // @[LoadQueue.scala 152:41:@13531.4]
  assign _T_15542 = addrQ_15 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@13532.4]
  assign conflict_15_7 = _T_15541 & _T_15542; // @[LoadQueue.scala 152:68:@13533.4]
  assign _T_15544 = entriesToCheck_15_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@13535.4]
  assign _T_15545 = _T_15544 & addrKnown_15; // @[LoadQueue.scala 152:41:@13536.4]
  assign _T_15546 = addrQ_15 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@13537.4]
  assign conflict_15_8 = _T_15545 & _T_15546; // @[LoadQueue.scala 152:68:@13538.4]
  assign _T_15548 = entriesToCheck_15_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@13540.4]
  assign _T_15549 = _T_15548 & addrKnown_15; // @[LoadQueue.scala 152:41:@13541.4]
  assign _T_15550 = addrQ_15 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@13542.4]
  assign conflict_15_9 = _T_15549 & _T_15550; // @[LoadQueue.scala 152:68:@13543.4]
  assign _T_15552 = entriesToCheck_15_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@13545.4]
  assign _T_15553 = _T_15552 & addrKnown_15; // @[LoadQueue.scala 152:41:@13546.4]
  assign _T_15554 = addrQ_15 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@13547.4]
  assign conflict_15_10 = _T_15553 & _T_15554; // @[LoadQueue.scala 152:68:@13548.4]
  assign _T_15556 = entriesToCheck_15_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@13550.4]
  assign _T_15557 = _T_15556 & addrKnown_15; // @[LoadQueue.scala 152:41:@13551.4]
  assign _T_15558 = addrQ_15 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@13552.4]
  assign conflict_15_11 = _T_15557 & _T_15558; // @[LoadQueue.scala 152:68:@13553.4]
  assign _T_15560 = entriesToCheck_15_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@13555.4]
  assign _T_15561 = _T_15560 & addrKnown_15; // @[LoadQueue.scala 152:41:@13556.4]
  assign _T_15562 = addrQ_15 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@13557.4]
  assign conflict_15_12 = _T_15561 & _T_15562; // @[LoadQueue.scala 152:68:@13558.4]
  assign _T_15564 = entriesToCheck_15_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@13560.4]
  assign _T_15565 = _T_15564 & addrKnown_15; // @[LoadQueue.scala 152:41:@13561.4]
  assign _T_15566 = addrQ_15 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@13562.4]
  assign conflict_15_13 = _T_15565 & _T_15566; // @[LoadQueue.scala 152:68:@13563.4]
  assign _T_15568 = entriesToCheck_15_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@13565.4]
  assign _T_15569 = _T_15568 & addrKnown_15; // @[LoadQueue.scala 152:41:@13566.4]
  assign _T_15570 = addrQ_15 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@13567.4]
  assign conflict_15_14 = _T_15569 & _T_15570; // @[LoadQueue.scala 152:68:@13568.4]
  assign _T_15572 = entriesToCheck_15_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@13570.4]
  assign _T_15573 = _T_15572 & addrKnown_15; // @[LoadQueue.scala 152:41:@13571.4]
  assign _T_15574 = addrQ_15 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@13572.4]
  assign conflict_15_15 = _T_15573 & _T_15574; // @[LoadQueue.scala 152:68:@13573.4]
  assign _T_16807 = io_storeAddrDone_0 == 1'h0; // @[LoadQueue.scala 163:13:@13576.4]
  assign storeAddrNotKnownFlags_0_0 = _T_16807 & entriesToCheck_0_0; // @[LoadQueue.scala 163:19:@13577.4]
  assign _T_16810 = io_storeAddrDone_1 == 1'h0; // @[LoadQueue.scala 163:13:@13578.4]
  assign storeAddrNotKnownFlags_0_1 = _T_16810 & entriesToCheck_0_1; // @[LoadQueue.scala 163:19:@13579.4]
  assign _T_16813 = io_storeAddrDone_2 == 1'h0; // @[LoadQueue.scala 163:13:@13580.4]
  assign storeAddrNotKnownFlags_0_2 = _T_16813 & entriesToCheck_0_2; // @[LoadQueue.scala 163:19:@13581.4]
  assign _T_16816 = io_storeAddrDone_3 == 1'h0; // @[LoadQueue.scala 163:13:@13582.4]
  assign storeAddrNotKnownFlags_0_3 = _T_16816 & entriesToCheck_0_3; // @[LoadQueue.scala 163:19:@13583.4]
  assign _T_16819 = io_storeAddrDone_4 == 1'h0; // @[LoadQueue.scala 163:13:@13584.4]
  assign storeAddrNotKnownFlags_0_4 = _T_16819 & entriesToCheck_0_4; // @[LoadQueue.scala 163:19:@13585.4]
  assign _T_16822 = io_storeAddrDone_5 == 1'h0; // @[LoadQueue.scala 163:13:@13586.4]
  assign storeAddrNotKnownFlags_0_5 = _T_16822 & entriesToCheck_0_5; // @[LoadQueue.scala 163:19:@13587.4]
  assign _T_16825 = io_storeAddrDone_6 == 1'h0; // @[LoadQueue.scala 163:13:@13588.4]
  assign storeAddrNotKnownFlags_0_6 = _T_16825 & entriesToCheck_0_6; // @[LoadQueue.scala 163:19:@13589.4]
  assign _T_16828 = io_storeAddrDone_7 == 1'h0; // @[LoadQueue.scala 163:13:@13590.4]
  assign storeAddrNotKnownFlags_0_7 = _T_16828 & entriesToCheck_0_7; // @[LoadQueue.scala 163:19:@13591.4]
  assign _T_16831 = io_storeAddrDone_8 == 1'h0; // @[LoadQueue.scala 163:13:@13592.4]
  assign storeAddrNotKnownFlags_0_8 = _T_16831 & entriesToCheck_0_8; // @[LoadQueue.scala 163:19:@13593.4]
  assign _T_16834 = io_storeAddrDone_9 == 1'h0; // @[LoadQueue.scala 163:13:@13594.4]
  assign storeAddrNotKnownFlags_0_9 = _T_16834 & entriesToCheck_0_9; // @[LoadQueue.scala 163:19:@13595.4]
  assign _T_16837 = io_storeAddrDone_10 == 1'h0; // @[LoadQueue.scala 163:13:@13596.4]
  assign storeAddrNotKnownFlags_0_10 = _T_16837 & entriesToCheck_0_10; // @[LoadQueue.scala 163:19:@13597.4]
  assign _T_16840 = io_storeAddrDone_11 == 1'h0; // @[LoadQueue.scala 163:13:@13598.4]
  assign storeAddrNotKnownFlags_0_11 = _T_16840 & entriesToCheck_0_11; // @[LoadQueue.scala 163:19:@13599.4]
  assign _T_16843 = io_storeAddrDone_12 == 1'h0; // @[LoadQueue.scala 163:13:@13600.4]
  assign storeAddrNotKnownFlags_0_12 = _T_16843 & entriesToCheck_0_12; // @[LoadQueue.scala 163:19:@13601.4]
  assign _T_16846 = io_storeAddrDone_13 == 1'h0; // @[LoadQueue.scala 163:13:@13602.4]
  assign storeAddrNotKnownFlags_0_13 = _T_16846 & entriesToCheck_0_13; // @[LoadQueue.scala 163:19:@13603.4]
  assign _T_16849 = io_storeAddrDone_14 == 1'h0; // @[LoadQueue.scala 163:13:@13604.4]
  assign storeAddrNotKnownFlags_0_14 = _T_16849 & entriesToCheck_0_14; // @[LoadQueue.scala 163:19:@13605.4]
  assign _T_16852 = io_storeAddrDone_15 == 1'h0; // @[LoadQueue.scala 163:13:@13606.4]
  assign storeAddrNotKnownFlags_0_15 = _T_16852 & entriesToCheck_0_15; // @[LoadQueue.scala 163:19:@13607.4]
  assign storeAddrNotKnownFlags_1_0 = _T_16807 & entriesToCheck_1_0; // @[LoadQueue.scala 163:19:@13625.4]
  assign storeAddrNotKnownFlags_1_1 = _T_16810 & entriesToCheck_1_1; // @[LoadQueue.scala 163:19:@13627.4]
  assign storeAddrNotKnownFlags_1_2 = _T_16813 & entriesToCheck_1_2; // @[LoadQueue.scala 163:19:@13629.4]
  assign storeAddrNotKnownFlags_1_3 = _T_16816 & entriesToCheck_1_3; // @[LoadQueue.scala 163:19:@13631.4]
  assign storeAddrNotKnownFlags_1_4 = _T_16819 & entriesToCheck_1_4; // @[LoadQueue.scala 163:19:@13633.4]
  assign storeAddrNotKnownFlags_1_5 = _T_16822 & entriesToCheck_1_5; // @[LoadQueue.scala 163:19:@13635.4]
  assign storeAddrNotKnownFlags_1_6 = _T_16825 & entriesToCheck_1_6; // @[LoadQueue.scala 163:19:@13637.4]
  assign storeAddrNotKnownFlags_1_7 = _T_16828 & entriesToCheck_1_7; // @[LoadQueue.scala 163:19:@13639.4]
  assign storeAddrNotKnownFlags_1_8 = _T_16831 & entriesToCheck_1_8; // @[LoadQueue.scala 163:19:@13641.4]
  assign storeAddrNotKnownFlags_1_9 = _T_16834 & entriesToCheck_1_9; // @[LoadQueue.scala 163:19:@13643.4]
  assign storeAddrNotKnownFlags_1_10 = _T_16837 & entriesToCheck_1_10; // @[LoadQueue.scala 163:19:@13645.4]
  assign storeAddrNotKnownFlags_1_11 = _T_16840 & entriesToCheck_1_11; // @[LoadQueue.scala 163:19:@13647.4]
  assign storeAddrNotKnownFlags_1_12 = _T_16843 & entriesToCheck_1_12; // @[LoadQueue.scala 163:19:@13649.4]
  assign storeAddrNotKnownFlags_1_13 = _T_16846 & entriesToCheck_1_13; // @[LoadQueue.scala 163:19:@13651.4]
  assign storeAddrNotKnownFlags_1_14 = _T_16849 & entriesToCheck_1_14; // @[LoadQueue.scala 163:19:@13653.4]
  assign storeAddrNotKnownFlags_1_15 = _T_16852 & entriesToCheck_1_15; // @[LoadQueue.scala 163:19:@13655.4]
  assign storeAddrNotKnownFlags_2_0 = _T_16807 & entriesToCheck_2_0; // @[LoadQueue.scala 163:19:@13673.4]
  assign storeAddrNotKnownFlags_2_1 = _T_16810 & entriesToCheck_2_1; // @[LoadQueue.scala 163:19:@13675.4]
  assign storeAddrNotKnownFlags_2_2 = _T_16813 & entriesToCheck_2_2; // @[LoadQueue.scala 163:19:@13677.4]
  assign storeAddrNotKnownFlags_2_3 = _T_16816 & entriesToCheck_2_3; // @[LoadQueue.scala 163:19:@13679.4]
  assign storeAddrNotKnownFlags_2_4 = _T_16819 & entriesToCheck_2_4; // @[LoadQueue.scala 163:19:@13681.4]
  assign storeAddrNotKnownFlags_2_5 = _T_16822 & entriesToCheck_2_5; // @[LoadQueue.scala 163:19:@13683.4]
  assign storeAddrNotKnownFlags_2_6 = _T_16825 & entriesToCheck_2_6; // @[LoadQueue.scala 163:19:@13685.4]
  assign storeAddrNotKnownFlags_2_7 = _T_16828 & entriesToCheck_2_7; // @[LoadQueue.scala 163:19:@13687.4]
  assign storeAddrNotKnownFlags_2_8 = _T_16831 & entriesToCheck_2_8; // @[LoadQueue.scala 163:19:@13689.4]
  assign storeAddrNotKnownFlags_2_9 = _T_16834 & entriesToCheck_2_9; // @[LoadQueue.scala 163:19:@13691.4]
  assign storeAddrNotKnownFlags_2_10 = _T_16837 & entriesToCheck_2_10; // @[LoadQueue.scala 163:19:@13693.4]
  assign storeAddrNotKnownFlags_2_11 = _T_16840 & entriesToCheck_2_11; // @[LoadQueue.scala 163:19:@13695.4]
  assign storeAddrNotKnownFlags_2_12 = _T_16843 & entriesToCheck_2_12; // @[LoadQueue.scala 163:19:@13697.4]
  assign storeAddrNotKnownFlags_2_13 = _T_16846 & entriesToCheck_2_13; // @[LoadQueue.scala 163:19:@13699.4]
  assign storeAddrNotKnownFlags_2_14 = _T_16849 & entriesToCheck_2_14; // @[LoadQueue.scala 163:19:@13701.4]
  assign storeAddrNotKnownFlags_2_15 = _T_16852 & entriesToCheck_2_15; // @[LoadQueue.scala 163:19:@13703.4]
  assign storeAddrNotKnownFlags_3_0 = _T_16807 & entriesToCheck_3_0; // @[LoadQueue.scala 163:19:@13721.4]
  assign storeAddrNotKnownFlags_3_1 = _T_16810 & entriesToCheck_3_1; // @[LoadQueue.scala 163:19:@13723.4]
  assign storeAddrNotKnownFlags_3_2 = _T_16813 & entriesToCheck_3_2; // @[LoadQueue.scala 163:19:@13725.4]
  assign storeAddrNotKnownFlags_3_3 = _T_16816 & entriesToCheck_3_3; // @[LoadQueue.scala 163:19:@13727.4]
  assign storeAddrNotKnownFlags_3_4 = _T_16819 & entriesToCheck_3_4; // @[LoadQueue.scala 163:19:@13729.4]
  assign storeAddrNotKnownFlags_3_5 = _T_16822 & entriesToCheck_3_5; // @[LoadQueue.scala 163:19:@13731.4]
  assign storeAddrNotKnownFlags_3_6 = _T_16825 & entriesToCheck_3_6; // @[LoadQueue.scala 163:19:@13733.4]
  assign storeAddrNotKnownFlags_3_7 = _T_16828 & entriesToCheck_3_7; // @[LoadQueue.scala 163:19:@13735.4]
  assign storeAddrNotKnownFlags_3_8 = _T_16831 & entriesToCheck_3_8; // @[LoadQueue.scala 163:19:@13737.4]
  assign storeAddrNotKnownFlags_3_9 = _T_16834 & entriesToCheck_3_9; // @[LoadQueue.scala 163:19:@13739.4]
  assign storeAddrNotKnownFlags_3_10 = _T_16837 & entriesToCheck_3_10; // @[LoadQueue.scala 163:19:@13741.4]
  assign storeAddrNotKnownFlags_3_11 = _T_16840 & entriesToCheck_3_11; // @[LoadQueue.scala 163:19:@13743.4]
  assign storeAddrNotKnownFlags_3_12 = _T_16843 & entriesToCheck_3_12; // @[LoadQueue.scala 163:19:@13745.4]
  assign storeAddrNotKnownFlags_3_13 = _T_16846 & entriesToCheck_3_13; // @[LoadQueue.scala 163:19:@13747.4]
  assign storeAddrNotKnownFlags_3_14 = _T_16849 & entriesToCheck_3_14; // @[LoadQueue.scala 163:19:@13749.4]
  assign storeAddrNotKnownFlags_3_15 = _T_16852 & entriesToCheck_3_15; // @[LoadQueue.scala 163:19:@13751.4]
  assign storeAddrNotKnownFlags_4_0 = _T_16807 & entriesToCheck_4_0; // @[LoadQueue.scala 163:19:@13769.4]
  assign storeAddrNotKnownFlags_4_1 = _T_16810 & entriesToCheck_4_1; // @[LoadQueue.scala 163:19:@13771.4]
  assign storeAddrNotKnownFlags_4_2 = _T_16813 & entriesToCheck_4_2; // @[LoadQueue.scala 163:19:@13773.4]
  assign storeAddrNotKnownFlags_4_3 = _T_16816 & entriesToCheck_4_3; // @[LoadQueue.scala 163:19:@13775.4]
  assign storeAddrNotKnownFlags_4_4 = _T_16819 & entriesToCheck_4_4; // @[LoadQueue.scala 163:19:@13777.4]
  assign storeAddrNotKnownFlags_4_5 = _T_16822 & entriesToCheck_4_5; // @[LoadQueue.scala 163:19:@13779.4]
  assign storeAddrNotKnownFlags_4_6 = _T_16825 & entriesToCheck_4_6; // @[LoadQueue.scala 163:19:@13781.4]
  assign storeAddrNotKnownFlags_4_7 = _T_16828 & entriesToCheck_4_7; // @[LoadQueue.scala 163:19:@13783.4]
  assign storeAddrNotKnownFlags_4_8 = _T_16831 & entriesToCheck_4_8; // @[LoadQueue.scala 163:19:@13785.4]
  assign storeAddrNotKnownFlags_4_9 = _T_16834 & entriesToCheck_4_9; // @[LoadQueue.scala 163:19:@13787.4]
  assign storeAddrNotKnownFlags_4_10 = _T_16837 & entriesToCheck_4_10; // @[LoadQueue.scala 163:19:@13789.4]
  assign storeAddrNotKnownFlags_4_11 = _T_16840 & entriesToCheck_4_11; // @[LoadQueue.scala 163:19:@13791.4]
  assign storeAddrNotKnownFlags_4_12 = _T_16843 & entriesToCheck_4_12; // @[LoadQueue.scala 163:19:@13793.4]
  assign storeAddrNotKnownFlags_4_13 = _T_16846 & entriesToCheck_4_13; // @[LoadQueue.scala 163:19:@13795.4]
  assign storeAddrNotKnownFlags_4_14 = _T_16849 & entriesToCheck_4_14; // @[LoadQueue.scala 163:19:@13797.4]
  assign storeAddrNotKnownFlags_4_15 = _T_16852 & entriesToCheck_4_15; // @[LoadQueue.scala 163:19:@13799.4]
  assign storeAddrNotKnownFlags_5_0 = _T_16807 & entriesToCheck_5_0; // @[LoadQueue.scala 163:19:@13817.4]
  assign storeAddrNotKnownFlags_5_1 = _T_16810 & entriesToCheck_5_1; // @[LoadQueue.scala 163:19:@13819.4]
  assign storeAddrNotKnownFlags_5_2 = _T_16813 & entriesToCheck_5_2; // @[LoadQueue.scala 163:19:@13821.4]
  assign storeAddrNotKnownFlags_5_3 = _T_16816 & entriesToCheck_5_3; // @[LoadQueue.scala 163:19:@13823.4]
  assign storeAddrNotKnownFlags_5_4 = _T_16819 & entriesToCheck_5_4; // @[LoadQueue.scala 163:19:@13825.4]
  assign storeAddrNotKnownFlags_5_5 = _T_16822 & entriesToCheck_5_5; // @[LoadQueue.scala 163:19:@13827.4]
  assign storeAddrNotKnownFlags_5_6 = _T_16825 & entriesToCheck_5_6; // @[LoadQueue.scala 163:19:@13829.4]
  assign storeAddrNotKnownFlags_5_7 = _T_16828 & entriesToCheck_5_7; // @[LoadQueue.scala 163:19:@13831.4]
  assign storeAddrNotKnownFlags_5_8 = _T_16831 & entriesToCheck_5_8; // @[LoadQueue.scala 163:19:@13833.4]
  assign storeAddrNotKnownFlags_5_9 = _T_16834 & entriesToCheck_5_9; // @[LoadQueue.scala 163:19:@13835.4]
  assign storeAddrNotKnownFlags_5_10 = _T_16837 & entriesToCheck_5_10; // @[LoadQueue.scala 163:19:@13837.4]
  assign storeAddrNotKnownFlags_5_11 = _T_16840 & entriesToCheck_5_11; // @[LoadQueue.scala 163:19:@13839.4]
  assign storeAddrNotKnownFlags_5_12 = _T_16843 & entriesToCheck_5_12; // @[LoadQueue.scala 163:19:@13841.4]
  assign storeAddrNotKnownFlags_5_13 = _T_16846 & entriesToCheck_5_13; // @[LoadQueue.scala 163:19:@13843.4]
  assign storeAddrNotKnownFlags_5_14 = _T_16849 & entriesToCheck_5_14; // @[LoadQueue.scala 163:19:@13845.4]
  assign storeAddrNotKnownFlags_5_15 = _T_16852 & entriesToCheck_5_15; // @[LoadQueue.scala 163:19:@13847.4]
  assign storeAddrNotKnownFlags_6_0 = _T_16807 & entriesToCheck_6_0; // @[LoadQueue.scala 163:19:@13865.4]
  assign storeAddrNotKnownFlags_6_1 = _T_16810 & entriesToCheck_6_1; // @[LoadQueue.scala 163:19:@13867.4]
  assign storeAddrNotKnownFlags_6_2 = _T_16813 & entriesToCheck_6_2; // @[LoadQueue.scala 163:19:@13869.4]
  assign storeAddrNotKnownFlags_6_3 = _T_16816 & entriesToCheck_6_3; // @[LoadQueue.scala 163:19:@13871.4]
  assign storeAddrNotKnownFlags_6_4 = _T_16819 & entriesToCheck_6_4; // @[LoadQueue.scala 163:19:@13873.4]
  assign storeAddrNotKnownFlags_6_5 = _T_16822 & entriesToCheck_6_5; // @[LoadQueue.scala 163:19:@13875.4]
  assign storeAddrNotKnownFlags_6_6 = _T_16825 & entriesToCheck_6_6; // @[LoadQueue.scala 163:19:@13877.4]
  assign storeAddrNotKnownFlags_6_7 = _T_16828 & entriesToCheck_6_7; // @[LoadQueue.scala 163:19:@13879.4]
  assign storeAddrNotKnownFlags_6_8 = _T_16831 & entriesToCheck_6_8; // @[LoadQueue.scala 163:19:@13881.4]
  assign storeAddrNotKnownFlags_6_9 = _T_16834 & entriesToCheck_6_9; // @[LoadQueue.scala 163:19:@13883.4]
  assign storeAddrNotKnownFlags_6_10 = _T_16837 & entriesToCheck_6_10; // @[LoadQueue.scala 163:19:@13885.4]
  assign storeAddrNotKnownFlags_6_11 = _T_16840 & entriesToCheck_6_11; // @[LoadQueue.scala 163:19:@13887.4]
  assign storeAddrNotKnownFlags_6_12 = _T_16843 & entriesToCheck_6_12; // @[LoadQueue.scala 163:19:@13889.4]
  assign storeAddrNotKnownFlags_6_13 = _T_16846 & entriesToCheck_6_13; // @[LoadQueue.scala 163:19:@13891.4]
  assign storeAddrNotKnownFlags_6_14 = _T_16849 & entriesToCheck_6_14; // @[LoadQueue.scala 163:19:@13893.4]
  assign storeAddrNotKnownFlags_6_15 = _T_16852 & entriesToCheck_6_15; // @[LoadQueue.scala 163:19:@13895.4]
  assign storeAddrNotKnownFlags_7_0 = _T_16807 & entriesToCheck_7_0; // @[LoadQueue.scala 163:19:@13913.4]
  assign storeAddrNotKnownFlags_7_1 = _T_16810 & entriesToCheck_7_1; // @[LoadQueue.scala 163:19:@13915.4]
  assign storeAddrNotKnownFlags_7_2 = _T_16813 & entriesToCheck_7_2; // @[LoadQueue.scala 163:19:@13917.4]
  assign storeAddrNotKnownFlags_7_3 = _T_16816 & entriesToCheck_7_3; // @[LoadQueue.scala 163:19:@13919.4]
  assign storeAddrNotKnownFlags_7_4 = _T_16819 & entriesToCheck_7_4; // @[LoadQueue.scala 163:19:@13921.4]
  assign storeAddrNotKnownFlags_7_5 = _T_16822 & entriesToCheck_7_5; // @[LoadQueue.scala 163:19:@13923.4]
  assign storeAddrNotKnownFlags_7_6 = _T_16825 & entriesToCheck_7_6; // @[LoadQueue.scala 163:19:@13925.4]
  assign storeAddrNotKnownFlags_7_7 = _T_16828 & entriesToCheck_7_7; // @[LoadQueue.scala 163:19:@13927.4]
  assign storeAddrNotKnownFlags_7_8 = _T_16831 & entriesToCheck_7_8; // @[LoadQueue.scala 163:19:@13929.4]
  assign storeAddrNotKnownFlags_7_9 = _T_16834 & entriesToCheck_7_9; // @[LoadQueue.scala 163:19:@13931.4]
  assign storeAddrNotKnownFlags_7_10 = _T_16837 & entriesToCheck_7_10; // @[LoadQueue.scala 163:19:@13933.4]
  assign storeAddrNotKnownFlags_7_11 = _T_16840 & entriesToCheck_7_11; // @[LoadQueue.scala 163:19:@13935.4]
  assign storeAddrNotKnownFlags_7_12 = _T_16843 & entriesToCheck_7_12; // @[LoadQueue.scala 163:19:@13937.4]
  assign storeAddrNotKnownFlags_7_13 = _T_16846 & entriesToCheck_7_13; // @[LoadQueue.scala 163:19:@13939.4]
  assign storeAddrNotKnownFlags_7_14 = _T_16849 & entriesToCheck_7_14; // @[LoadQueue.scala 163:19:@13941.4]
  assign storeAddrNotKnownFlags_7_15 = _T_16852 & entriesToCheck_7_15; // @[LoadQueue.scala 163:19:@13943.4]
  assign storeAddrNotKnownFlags_8_0 = _T_16807 & entriesToCheck_8_0; // @[LoadQueue.scala 163:19:@13961.4]
  assign storeAddrNotKnownFlags_8_1 = _T_16810 & entriesToCheck_8_1; // @[LoadQueue.scala 163:19:@13963.4]
  assign storeAddrNotKnownFlags_8_2 = _T_16813 & entriesToCheck_8_2; // @[LoadQueue.scala 163:19:@13965.4]
  assign storeAddrNotKnownFlags_8_3 = _T_16816 & entriesToCheck_8_3; // @[LoadQueue.scala 163:19:@13967.4]
  assign storeAddrNotKnownFlags_8_4 = _T_16819 & entriesToCheck_8_4; // @[LoadQueue.scala 163:19:@13969.4]
  assign storeAddrNotKnownFlags_8_5 = _T_16822 & entriesToCheck_8_5; // @[LoadQueue.scala 163:19:@13971.4]
  assign storeAddrNotKnownFlags_8_6 = _T_16825 & entriesToCheck_8_6; // @[LoadQueue.scala 163:19:@13973.4]
  assign storeAddrNotKnownFlags_8_7 = _T_16828 & entriesToCheck_8_7; // @[LoadQueue.scala 163:19:@13975.4]
  assign storeAddrNotKnownFlags_8_8 = _T_16831 & entriesToCheck_8_8; // @[LoadQueue.scala 163:19:@13977.4]
  assign storeAddrNotKnownFlags_8_9 = _T_16834 & entriesToCheck_8_9; // @[LoadQueue.scala 163:19:@13979.4]
  assign storeAddrNotKnownFlags_8_10 = _T_16837 & entriesToCheck_8_10; // @[LoadQueue.scala 163:19:@13981.4]
  assign storeAddrNotKnownFlags_8_11 = _T_16840 & entriesToCheck_8_11; // @[LoadQueue.scala 163:19:@13983.4]
  assign storeAddrNotKnownFlags_8_12 = _T_16843 & entriesToCheck_8_12; // @[LoadQueue.scala 163:19:@13985.4]
  assign storeAddrNotKnownFlags_8_13 = _T_16846 & entriesToCheck_8_13; // @[LoadQueue.scala 163:19:@13987.4]
  assign storeAddrNotKnownFlags_8_14 = _T_16849 & entriesToCheck_8_14; // @[LoadQueue.scala 163:19:@13989.4]
  assign storeAddrNotKnownFlags_8_15 = _T_16852 & entriesToCheck_8_15; // @[LoadQueue.scala 163:19:@13991.4]
  assign storeAddrNotKnownFlags_9_0 = _T_16807 & entriesToCheck_9_0; // @[LoadQueue.scala 163:19:@14009.4]
  assign storeAddrNotKnownFlags_9_1 = _T_16810 & entriesToCheck_9_1; // @[LoadQueue.scala 163:19:@14011.4]
  assign storeAddrNotKnownFlags_9_2 = _T_16813 & entriesToCheck_9_2; // @[LoadQueue.scala 163:19:@14013.4]
  assign storeAddrNotKnownFlags_9_3 = _T_16816 & entriesToCheck_9_3; // @[LoadQueue.scala 163:19:@14015.4]
  assign storeAddrNotKnownFlags_9_4 = _T_16819 & entriesToCheck_9_4; // @[LoadQueue.scala 163:19:@14017.4]
  assign storeAddrNotKnownFlags_9_5 = _T_16822 & entriesToCheck_9_5; // @[LoadQueue.scala 163:19:@14019.4]
  assign storeAddrNotKnownFlags_9_6 = _T_16825 & entriesToCheck_9_6; // @[LoadQueue.scala 163:19:@14021.4]
  assign storeAddrNotKnownFlags_9_7 = _T_16828 & entriesToCheck_9_7; // @[LoadQueue.scala 163:19:@14023.4]
  assign storeAddrNotKnownFlags_9_8 = _T_16831 & entriesToCheck_9_8; // @[LoadQueue.scala 163:19:@14025.4]
  assign storeAddrNotKnownFlags_9_9 = _T_16834 & entriesToCheck_9_9; // @[LoadQueue.scala 163:19:@14027.4]
  assign storeAddrNotKnownFlags_9_10 = _T_16837 & entriesToCheck_9_10; // @[LoadQueue.scala 163:19:@14029.4]
  assign storeAddrNotKnownFlags_9_11 = _T_16840 & entriesToCheck_9_11; // @[LoadQueue.scala 163:19:@14031.4]
  assign storeAddrNotKnownFlags_9_12 = _T_16843 & entriesToCheck_9_12; // @[LoadQueue.scala 163:19:@14033.4]
  assign storeAddrNotKnownFlags_9_13 = _T_16846 & entriesToCheck_9_13; // @[LoadQueue.scala 163:19:@14035.4]
  assign storeAddrNotKnownFlags_9_14 = _T_16849 & entriesToCheck_9_14; // @[LoadQueue.scala 163:19:@14037.4]
  assign storeAddrNotKnownFlags_9_15 = _T_16852 & entriesToCheck_9_15; // @[LoadQueue.scala 163:19:@14039.4]
  assign storeAddrNotKnownFlags_10_0 = _T_16807 & entriesToCheck_10_0; // @[LoadQueue.scala 163:19:@14057.4]
  assign storeAddrNotKnownFlags_10_1 = _T_16810 & entriesToCheck_10_1; // @[LoadQueue.scala 163:19:@14059.4]
  assign storeAddrNotKnownFlags_10_2 = _T_16813 & entriesToCheck_10_2; // @[LoadQueue.scala 163:19:@14061.4]
  assign storeAddrNotKnownFlags_10_3 = _T_16816 & entriesToCheck_10_3; // @[LoadQueue.scala 163:19:@14063.4]
  assign storeAddrNotKnownFlags_10_4 = _T_16819 & entriesToCheck_10_4; // @[LoadQueue.scala 163:19:@14065.4]
  assign storeAddrNotKnownFlags_10_5 = _T_16822 & entriesToCheck_10_5; // @[LoadQueue.scala 163:19:@14067.4]
  assign storeAddrNotKnownFlags_10_6 = _T_16825 & entriesToCheck_10_6; // @[LoadQueue.scala 163:19:@14069.4]
  assign storeAddrNotKnownFlags_10_7 = _T_16828 & entriesToCheck_10_7; // @[LoadQueue.scala 163:19:@14071.4]
  assign storeAddrNotKnownFlags_10_8 = _T_16831 & entriesToCheck_10_8; // @[LoadQueue.scala 163:19:@14073.4]
  assign storeAddrNotKnownFlags_10_9 = _T_16834 & entriesToCheck_10_9; // @[LoadQueue.scala 163:19:@14075.4]
  assign storeAddrNotKnownFlags_10_10 = _T_16837 & entriesToCheck_10_10; // @[LoadQueue.scala 163:19:@14077.4]
  assign storeAddrNotKnownFlags_10_11 = _T_16840 & entriesToCheck_10_11; // @[LoadQueue.scala 163:19:@14079.4]
  assign storeAddrNotKnownFlags_10_12 = _T_16843 & entriesToCheck_10_12; // @[LoadQueue.scala 163:19:@14081.4]
  assign storeAddrNotKnownFlags_10_13 = _T_16846 & entriesToCheck_10_13; // @[LoadQueue.scala 163:19:@14083.4]
  assign storeAddrNotKnownFlags_10_14 = _T_16849 & entriesToCheck_10_14; // @[LoadQueue.scala 163:19:@14085.4]
  assign storeAddrNotKnownFlags_10_15 = _T_16852 & entriesToCheck_10_15; // @[LoadQueue.scala 163:19:@14087.4]
  assign storeAddrNotKnownFlags_11_0 = _T_16807 & entriesToCheck_11_0; // @[LoadQueue.scala 163:19:@14105.4]
  assign storeAddrNotKnownFlags_11_1 = _T_16810 & entriesToCheck_11_1; // @[LoadQueue.scala 163:19:@14107.4]
  assign storeAddrNotKnownFlags_11_2 = _T_16813 & entriesToCheck_11_2; // @[LoadQueue.scala 163:19:@14109.4]
  assign storeAddrNotKnownFlags_11_3 = _T_16816 & entriesToCheck_11_3; // @[LoadQueue.scala 163:19:@14111.4]
  assign storeAddrNotKnownFlags_11_4 = _T_16819 & entriesToCheck_11_4; // @[LoadQueue.scala 163:19:@14113.4]
  assign storeAddrNotKnownFlags_11_5 = _T_16822 & entriesToCheck_11_5; // @[LoadQueue.scala 163:19:@14115.4]
  assign storeAddrNotKnownFlags_11_6 = _T_16825 & entriesToCheck_11_6; // @[LoadQueue.scala 163:19:@14117.4]
  assign storeAddrNotKnownFlags_11_7 = _T_16828 & entriesToCheck_11_7; // @[LoadQueue.scala 163:19:@14119.4]
  assign storeAddrNotKnownFlags_11_8 = _T_16831 & entriesToCheck_11_8; // @[LoadQueue.scala 163:19:@14121.4]
  assign storeAddrNotKnownFlags_11_9 = _T_16834 & entriesToCheck_11_9; // @[LoadQueue.scala 163:19:@14123.4]
  assign storeAddrNotKnownFlags_11_10 = _T_16837 & entriesToCheck_11_10; // @[LoadQueue.scala 163:19:@14125.4]
  assign storeAddrNotKnownFlags_11_11 = _T_16840 & entriesToCheck_11_11; // @[LoadQueue.scala 163:19:@14127.4]
  assign storeAddrNotKnownFlags_11_12 = _T_16843 & entriesToCheck_11_12; // @[LoadQueue.scala 163:19:@14129.4]
  assign storeAddrNotKnownFlags_11_13 = _T_16846 & entriesToCheck_11_13; // @[LoadQueue.scala 163:19:@14131.4]
  assign storeAddrNotKnownFlags_11_14 = _T_16849 & entriesToCheck_11_14; // @[LoadQueue.scala 163:19:@14133.4]
  assign storeAddrNotKnownFlags_11_15 = _T_16852 & entriesToCheck_11_15; // @[LoadQueue.scala 163:19:@14135.4]
  assign storeAddrNotKnownFlags_12_0 = _T_16807 & entriesToCheck_12_0; // @[LoadQueue.scala 163:19:@14153.4]
  assign storeAddrNotKnownFlags_12_1 = _T_16810 & entriesToCheck_12_1; // @[LoadQueue.scala 163:19:@14155.4]
  assign storeAddrNotKnownFlags_12_2 = _T_16813 & entriesToCheck_12_2; // @[LoadQueue.scala 163:19:@14157.4]
  assign storeAddrNotKnownFlags_12_3 = _T_16816 & entriesToCheck_12_3; // @[LoadQueue.scala 163:19:@14159.4]
  assign storeAddrNotKnownFlags_12_4 = _T_16819 & entriesToCheck_12_4; // @[LoadQueue.scala 163:19:@14161.4]
  assign storeAddrNotKnownFlags_12_5 = _T_16822 & entriesToCheck_12_5; // @[LoadQueue.scala 163:19:@14163.4]
  assign storeAddrNotKnownFlags_12_6 = _T_16825 & entriesToCheck_12_6; // @[LoadQueue.scala 163:19:@14165.4]
  assign storeAddrNotKnownFlags_12_7 = _T_16828 & entriesToCheck_12_7; // @[LoadQueue.scala 163:19:@14167.4]
  assign storeAddrNotKnownFlags_12_8 = _T_16831 & entriesToCheck_12_8; // @[LoadQueue.scala 163:19:@14169.4]
  assign storeAddrNotKnownFlags_12_9 = _T_16834 & entriesToCheck_12_9; // @[LoadQueue.scala 163:19:@14171.4]
  assign storeAddrNotKnownFlags_12_10 = _T_16837 & entriesToCheck_12_10; // @[LoadQueue.scala 163:19:@14173.4]
  assign storeAddrNotKnownFlags_12_11 = _T_16840 & entriesToCheck_12_11; // @[LoadQueue.scala 163:19:@14175.4]
  assign storeAddrNotKnownFlags_12_12 = _T_16843 & entriesToCheck_12_12; // @[LoadQueue.scala 163:19:@14177.4]
  assign storeAddrNotKnownFlags_12_13 = _T_16846 & entriesToCheck_12_13; // @[LoadQueue.scala 163:19:@14179.4]
  assign storeAddrNotKnownFlags_12_14 = _T_16849 & entriesToCheck_12_14; // @[LoadQueue.scala 163:19:@14181.4]
  assign storeAddrNotKnownFlags_12_15 = _T_16852 & entriesToCheck_12_15; // @[LoadQueue.scala 163:19:@14183.4]
  assign storeAddrNotKnownFlags_13_0 = _T_16807 & entriesToCheck_13_0; // @[LoadQueue.scala 163:19:@14201.4]
  assign storeAddrNotKnownFlags_13_1 = _T_16810 & entriesToCheck_13_1; // @[LoadQueue.scala 163:19:@14203.4]
  assign storeAddrNotKnownFlags_13_2 = _T_16813 & entriesToCheck_13_2; // @[LoadQueue.scala 163:19:@14205.4]
  assign storeAddrNotKnownFlags_13_3 = _T_16816 & entriesToCheck_13_3; // @[LoadQueue.scala 163:19:@14207.4]
  assign storeAddrNotKnownFlags_13_4 = _T_16819 & entriesToCheck_13_4; // @[LoadQueue.scala 163:19:@14209.4]
  assign storeAddrNotKnownFlags_13_5 = _T_16822 & entriesToCheck_13_5; // @[LoadQueue.scala 163:19:@14211.4]
  assign storeAddrNotKnownFlags_13_6 = _T_16825 & entriesToCheck_13_6; // @[LoadQueue.scala 163:19:@14213.4]
  assign storeAddrNotKnownFlags_13_7 = _T_16828 & entriesToCheck_13_7; // @[LoadQueue.scala 163:19:@14215.4]
  assign storeAddrNotKnownFlags_13_8 = _T_16831 & entriesToCheck_13_8; // @[LoadQueue.scala 163:19:@14217.4]
  assign storeAddrNotKnownFlags_13_9 = _T_16834 & entriesToCheck_13_9; // @[LoadQueue.scala 163:19:@14219.4]
  assign storeAddrNotKnownFlags_13_10 = _T_16837 & entriesToCheck_13_10; // @[LoadQueue.scala 163:19:@14221.4]
  assign storeAddrNotKnownFlags_13_11 = _T_16840 & entriesToCheck_13_11; // @[LoadQueue.scala 163:19:@14223.4]
  assign storeAddrNotKnownFlags_13_12 = _T_16843 & entriesToCheck_13_12; // @[LoadQueue.scala 163:19:@14225.4]
  assign storeAddrNotKnownFlags_13_13 = _T_16846 & entriesToCheck_13_13; // @[LoadQueue.scala 163:19:@14227.4]
  assign storeAddrNotKnownFlags_13_14 = _T_16849 & entriesToCheck_13_14; // @[LoadQueue.scala 163:19:@14229.4]
  assign storeAddrNotKnownFlags_13_15 = _T_16852 & entriesToCheck_13_15; // @[LoadQueue.scala 163:19:@14231.4]
  assign storeAddrNotKnownFlags_14_0 = _T_16807 & entriesToCheck_14_0; // @[LoadQueue.scala 163:19:@14249.4]
  assign storeAddrNotKnownFlags_14_1 = _T_16810 & entriesToCheck_14_1; // @[LoadQueue.scala 163:19:@14251.4]
  assign storeAddrNotKnownFlags_14_2 = _T_16813 & entriesToCheck_14_2; // @[LoadQueue.scala 163:19:@14253.4]
  assign storeAddrNotKnownFlags_14_3 = _T_16816 & entriesToCheck_14_3; // @[LoadQueue.scala 163:19:@14255.4]
  assign storeAddrNotKnownFlags_14_4 = _T_16819 & entriesToCheck_14_4; // @[LoadQueue.scala 163:19:@14257.4]
  assign storeAddrNotKnownFlags_14_5 = _T_16822 & entriesToCheck_14_5; // @[LoadQueue.scala 163:19:@14259.4]
  assign storeAddrNotKnownFlags_14_6 = _T_16825 & entriesToCheck_14_6; // @[LoadQueue.scala 163:19:@14261.4]
  assign storeAddrNotKnownFlags_14_7 = _T_16828 & entriesToCheck_14_7; // @[LoadQueue.scala 163:19:@14263.4]
  assign storeAddrNotKnownFlags_14_8 = _T_16831 & entriesToCheck_14_8; // @[LoadQueue.scala 163:19:@14265.4]
  assign storeAddrNotKnownFlags_14_9 = _T_16834 & entriesToCheck_14_9; // @[LoadQueue.scala 163:19:@14267.4]
  assign storeAddrNotKnownFlags_14_10 = _T_16837 & entriesToCheck_14_10; // @[LoadQueue.scala 163:19:@14269.4]
  assign storeAddrNotKnownFlags_14_11 = _T_16840 & entriesToCheck_14_11; // @[LoadQueue.scala 163:19:@14271.4]
  assign storeAddrNotKnownFlags_14_12 = _T_16843 & entriesToCheck_14_12; // @[LoadQueue.scala 163:19:@14273.4]
  assign storeAddrNotKnownFlags_14_13 = _T_16846 & entriesToCheck_14_13; // @[LoadQueue.scala 163:19:@14275.4]
  assign storeAddrNotKnownFlags_14_14 = _T_16849 & entriesToCheck_14_14; // @[LoadQueue.scala 163:19:@14277.4]
  assign storeAddrNotKnownFlags_14_15 = _T_16852 & entriesToCheck_14_15; // @[LoadQueue.scala 163:19:@14279.4]
  assign storeAddrNotKnownFlags_15_0 = _T_16807 & entriesToCheck_15_0; // @[LoadQueue.scala 163:19:@14297.4]
  assign storeAddrNotKnownFlags_15_1 = _T_16810 & entriesToCheck_15_1; // @[LoadQueue.scala 163:19:@14299.4]
  assign storeAddrNotKnownFlags_15_2 = _T_16813 & entriesToCheck_15_2; // @[LoadQueue.scala 163:19:@14301.4]
  assign storeAddrNotKnownFlags_15_3 = _T_16816 & entriesToCheck_15_3; // @[LoadQueue.scala 163:19:@14303.4]
  assign storeAddrNotKnownFlags_15_4 = _T_16819 & entriesToCheck_15_4; // @[LoadQueue.scala 163:19:@14305.4]
  assign storeAddrNotKnownFlags_15_5 = _T_16822 & entriesToCheck_15_5; // @[LoadQueue.scala 163:19:@14307.4]
  assign storeAddrNotKnownFlags_15_6 = _T_16825 & entriesToCheck_15_6; // @[LoadQueue.scala 163:19:@14309.4]
  assign storeAddrNotKnownFlags_15_7 = _T_16828 & entriesToCheck_15_7; // @[LoadQueue.scala 163:19:@14311.4]
  assign storeAddrNotKnownFlags_15_8 = _T_16831 & entriesToCheck_15_8; // @[LoadQueue.scala 163:19:@14313.4]
  assign storeAddrNotKnownFlags_15_9 = _T_16834 & entriesToCheck_15_9; // @[LoadQueue.scala 163:19:@14315.4]
  assign storeAddrNotKnownFlags_15_10 = _T_16837 & entriesToCheck_15_10; // @[LoadQueue.scala 163:19:@14317.4]
  assign storeAddrNotKnownFlags_15_11 = _T_16840 & entriesToCheck_15_11; // @[LoadQueue.scala 163:19:@14319.4]
  assign storeAddrNotKnownFlags_15_12 = _T_16843 & entriesToCheck_15_12; // @[LoadQueue.scala 163:19:@14321.4]
  assign storeAddrNotKnownFlags_15_13 = _T_16846 & entriesToCheck_15_13; // @[LoadQueue.scala 163:19:@14323.4]
  assign storeAddrNotKnownFlags_15_14 = _T_16849 & entriesToCheck_15_14; // @[LoadQueue.scala 163:19:@14325.4]
  assign storeAddrNotKnownFlags_15_15 = _T_16852 & entriesToCheck_15_15; // @[LoadQueue.scala 163:19:@14327.4]
  assign _T_18010 = {conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0}; // @[Mux.scala 19:72:@14658.4]
  assign _T_18017 = {conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8}; // @[Mux.scala 19:72:@14665.4]
  assign _T_18018 = {conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,_T_18010}; // @[Mux.scala 19:72:@14666.4]
  assign _T_18020 = _T_2697 ? _T_18018 : 16'h0; // @[Mux.scala 19:72:@14667.4]
  assign _T_18027 = {conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1}; // @[Mux.scala 19:72:@14674.4]
  assign _T_18034 = {conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9}; // @[Mux.scala 19:72:@14681.4]
  assign _T_18035 = {conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,_T_18027}; // @[Mux.scala 19:72:@14682.4]
  assign _T_18037 = _T_2698 ? _T_18035 : 16'h0; // @[Mux.scala 19:72:@14683.4]
  assign _T_18044 = {conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2}; // @[Mux.scala 19:72:@14690.4]
  assign _T_18051 = {conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10}; // @[Mux.scala 19:72:@14697.4]
  assign _T_18052 = {conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,_T_18044}; // @[Mux.scala 19:72:@14698.4]
  assign _T_18054 = _T_2699 ? _T_18052 : 16'h0; // @[Mux.scala 19:72:@14699.4]
  assign _T_18061 = {conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3}; // @[Mux.scala 19:72:@14706.4]
  assign _T_18068 = {conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11}; // @[Mux.scala 19:72:@14713.4]
  assign _T_18069 = {conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,_T_18061}; // @[Mux.scala 19:72:@14714.4]
  assign _T_18071 = _T_2700 ? _T_18069 : 16'h0; // @[Mux.scala 19:72:@14715.4]
  assign _T_18078 = {conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4}; // @[Mux.scala 19:72:@14722.4]
  assign _T_18085 = {conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12}; // @[Mux.scala 19:72:@14729.4]
  assign _T_18086 = {conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,_T_18078}; // @[Mux.scala 19:72:@14730.4]
  assign _T_18088 = _T_2701 ? _T_18086 : 16'h0; // @[Mux.scala 19:72:@14731.4]
  assign _T_18095 = {conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5}; // @[Mux.scala 19:72:@14738.4]
  assign _T_18102 = {conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13}; // @[Mux.scala 19:72:@14745.4]
  assign _T_18103 = {conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,_T_18095}; // @[Mux.scala 19:72:@14746.4]
  assign _T_18105 = _T_2702 ? _T_18103 : 16'h0; // @[Mux.scala 19:72:@14747.4]
  assign _T_18112 = {conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6}; // @[Mux.scala 19:72:@14754.4]
  assign _T_18119 = {conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14}; // @[Mux.scala 19:72:@14761.4]
  assign _T_18120 = {conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,_T_18112}; // @[Mux.scala 19:72:@14762.4]
  assign _T_18122 = _T_2703 ? _T_18120 : 16'h0; // @[Mux.scala 19:72:@14763.4]
  assign _T_18129 = {conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7}; // @[Mux.scala 19:72:@14770.4]
  assign _T_18136 = {conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15}; // @[Mux.scala 19:72:@14777.4]
  assign _T_18137 = {conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,_T_18129}; // @[Mux.scala 19:72:@14778.4]
  assign _T_18139 = _T_2704 ? _T_18137 : 16'h0; // @[Mux.scala 19:72:@14779.4]
  assign _T_18154 = {conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,_T_18017}; // @[Mux.scala 19:72:@14794.4]
  assign _T_18156 = _T_2705 ? _T_18154 : 16'h0; // @[Mux.scala 19:72:@14795.4]
  assign _T_18171 = {conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,_T_18034}; // @[Mux.scala 19:72:@14810.4]
  assign _T_18173 = _T_2706 ? _T_18171 : 16'h0; // @[Mux.scala 19:72:@14811.4]
  assign _T_18188 = {conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,_T_18051}; // @[Mux.scala 19:72:@14826.4]
  assign _T_18190 = _T_2707 ? _T_18188 : 16'h0; // @[Mux.scala 19:72:@14827.4]
  assign _T_18205 = {conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,_T_18068}; // @[Mux.scala 19:72:@14842.4]
  assign _T_18207 = _T_2708 ? _T_18205 : 16'h0; // @[Mux.scala 19:72:@14843.4]
  assign _T_18222 = {conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,_T_18085}; // @[Mux.scala 19:72:@14858.4]
  assign _T_18224 = _T_2709 ? _T_18222 : 16'h0; // @[Mux.scala 19:72:@14859.4]
  assign _T_18239 = {conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,_T_18102}; // @[Mux.scala 19:72:@14874.4]
  assign _T_18241 = _T_2710 ? _T_18239 : 16'h0; // @[Mux.scala 19:72:@14875.4]
  assign _T_18256 = {conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,_T_18119}; // @[Mux.scala 19:72:@14890.4]
  assign _T_18258 = _T_2711 ? _T_18256 : 16'h0; // @[Mux.scala 19:72:@14891.4]
  assign _T_18273 = {conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,_T_18136}; // @[Mux.scala 19:72:@14906.4]
  assign _T_18275 = _T_2712 ? _T_18273 : 16'h0; // @[Mux.scala 19:72:@14907.4]
  assign _T_18276 = _T_18020 | _T_18037; // @[Mux.scala 19:72:@14908.4]
  assign _T_18277 = _T_18276 | _T_18054; // @[Mux.scala 19:72:@14909.4]
  assign _T_18278 = _T_18277 | _T_18071; // @[Mux.scala 19:72:@14910.4]
  assign _T_18279 = _T_18278 | _T_18088; // @[Mux.scala 19:72:@14911.4]
  assign _T_18280 = _T_18279 | _T_18105; // @[Mux.scala 19:72:@14912.4]
  assign _T_18281 = _T_18280 | _T_18122; // @[Mux.scala 19:72:@14913.4]
  assign _T_18282 = _T_18281 | _T_18139; // @[Mux.scala 19:72:@14914.4]
  assign _T_18283 = _T_18282 | _T_18156; // @[Mux.scala 19:72:@14915.4]
  assign _T_18284 = _T_18283 | _T_18173; // @[Mux.scala 19:72:@14916.4]
  assign _T_18285 = _T_18284 | _T_18190; // @[Mux.scala 19:72:@14917.4]
  assign _T_18286 = _T_18285 | _T_18207; // @[Mux.scala 19:72:@14918.4]
  assign _T_18287 = _T_18286 | _T_18224; // @[Mux.scala 19:72:@14919.4]
  assign _T_18288 = _T_18287 | _T_18241; // @[Mux.scala 19:72:@14920.4]
  assign _T_18289 = _T_18288 | _T_18258; // @[Mux.scala 19:72:@14921.4]
  assign _T_18290 = _T_18289 | _T_18275; // @[Mux.scala 19:72:@14922.4]
  assign _T_18868 = {conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0}; // @[Mux.scala 19:72:@15272.4]
  assign _T_18875 = {conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8}; // @[Mux.scala 19:72:@15279.4]
  assign _T_18876 = {conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,_T_18868}; // @[Mux.scala 19:72:@15280.4]
  assign _T_18878 = _T_2697 ? _T_18876 : 16'h0; // @[Mux.scala 19:72:@15281.4]
  assign _T_18885 = {conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1}; // @[Mux.scala 19:72:@15288.4]
  assign _T_18892 = {conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9}; // @[Mux.scala 19:72:@15295.4]
  assign _T_18893 = {conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,_T_18885}; // @[Mux.scala 19:72:@15296.4]
  assign _T_18895 = _T_2698 ? _T_18893 : 16'h0; // @[Mux.scala 19:72:@15297.4]
  assign _T_18902 = {conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2}; // @[Mux.scala 19:72:@15304.4]
  assign _T_18909 = {conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10}; // @[Mux.scala 19:72:@15311.4]
  assign _T_18910 = {conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,_T_18902}; // @[Mux.scala 19:72:@15312.4]
  assign _T_18912 = _T_2699 ? _T_18910 : 16'h0; // @[Mux.scala 19:72:@15313.4]
  assign _T_18919 = {conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3}; // @[Mux.scala 19:72:@15320.4]
  assign _T_18926 = {conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11}; // @[Mux.scala 19:72:@15327.4]
  assign _T_18927 = {conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,_T_18919}; // @[Mux.scala 19:72:@15328.4]
  assign _T_18929 = _T_2700 ? _T_18927 : 16'h0; // @[Mux.scala 19:72:@15329.4]
  assign _T_18936 = {conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4}; // @[Mux.scala 19:72:@15336.4]
  assign _T_18943 = {conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12}; // @[Mux.scala 19:72:@15343.4]
  assign _T_18944 = {conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,_T_18936}; // @[Mux.scala 19:72:@15344.4]
  assign _T_18946 = _T_2701 ? _T_18944 : 16'h0; // @[Mux.scala 19:72:@15345.4]
  assign _T_18953 = {conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5}; // @[Mux.scala 19:72:@15352.4]
  assign _T_18960 = {conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13}; // @[Mux.scala 19:72:@15359.4]
  assign _T_18961 = {conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,_T_18953}; // @[Mux.scala 19:72:@15360.4]
  assign _T_18963 = _T_2702 ? _T_18961 : 16'h0; // @[Mux.scala 19:72:@15361.4]
  assign _T_18970 = {conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6}; // @[Mux.scala 19:72:@15368.4]
  assign _T_18977 = {conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14}; // @[Mux.scala 19:72:@15375.4]
  assign _T_18978 = {conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,_T_18970}; // @[Mux.scala 19:72:@15376.4]
  assign _T_18980 = _T_2703 ? _T_18978 : 16'h0; // @[Mux.scala 19:72:@15377.4]
  assign _T_18987 = {conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7}; // @[Mux.scala 19:72:@15384.4]
  assign _T_18994 = {conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15}; // @[Mux.scala 19:72:@15391.4]
  assign _T_18995 = {conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,_T_18987}; // @[Mux.scala 19:72:@15392.4]
  assign _T_18997 = _T_2704 ? _T_18995 : 16'h0; // @[Mux.scala 19:72:@15393.4]
  assign _T_19012 = {conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,_T_18875}; // @[Mux.scala 19:72:@15408.4]
  assign _T_19014 = _T_2705 ? _T_19012 : 16'h0; // @[Mux.scala 19:72:@15409.4]
  assign _T_19029 = {conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,_T_18892}; // @[Mux.scala 19:72:@15424.4]
  assign _T_19031 = _T_2706 ? _T_19029 : 16'h0; // @[Mux.scala 19:72:@15425.4]
  assign _T_19046 = {conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,_T_18909}; // @[Mux.scala 19:72:@15440.4]
  assign _T_19048 = _T_2707 ? _T_19046 : 16'h0; // @[Mux.scala 19:72:@15441.4]
  assign _T_19063 = {conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,_T_18926}; // @[Mux.scala 19:72:@15456.4]
  assign _T_19065 = _T_2708 ? _T_19063 : 16'h0; // @[Mux.scala 19:72:@15457.4]
  assign _T_19080 = {conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,_T_18943}; // @[Mux.scala 19:72:@15472.4]
  assign _T_19082 = _T_2709 ? _T_19080 : 16'h0; // @[Mux.scala 19:72:@15473.4]
  assign _T_19097 = {conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,_T_18960}; // @[Mux.scala 19:72:@15488.4]
  assign _T_19099 = _T_2710 ? _T_19097 : 16'h0; // @[Mux.scala 19:72:@15489.4]
  assign _T_19114 = {conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,_T_18977}; // @[Mux.scala 19:72:@15504.4]
  assign _T_19116 = _T_2711 ? _T_19114 : 16'h0; // @[Mux.scala 19:72:@15505.4]
  assign _T_19131 = {conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,_T_18994}; // @[Mux.scala 19:72:@15520.4]
  assign _T_19133 = _T_2712 ? _T_19131 : 16'h0; // @[Mux.scala 19:72:@15521.4]
  assign _T_19134 = _T_18878 | _T_18895; // @[Mux.scala 19:72:@15522.4]
  assign _T_19135 = _T_19134 | _T_18912; // @[Mux.scala 19:72:@15523.4]
  assign _T_19136 = _T_19135 | _T_18929; // @[Mux.scala 19:72:@15524.4]
  assign _T_19137 = _T_19136 | _T_18946; // @[Mux.scala 19:72:@15525.4]
  assign _T_19138 = _T_19137 | _T_18963; // @[Mux.scala 19:72:@15526.4]
  assign _T_19139 = _T_19138 | _T_18980; // @[Mux.scala 19:72:@15527.4]
  assign _T_19140 = _T_19139 | _T_18997; // @[Mux.scala 19:72:@15528.4]
  assign _T_19141 = _T_19140 | _T_19014; // @[Mux.scala 19:72:@15529.4]
  assign _T_19142 = _T_19141 | _T_19031; // @[Mux.scala 19:72:@15530.4]
  assign _T_19143 = _T_19142 | _T_19048; // @[Mux.scala 19:72:@15531.4]
  assign _T_19144 = _T_19143 | _T_19065; // @[Mux.scala 19:72:@15532.4]
  assign _T_19145 = _T_19144 | _T_19082; // @[Mux.scala 19:72:@15533.4]
  assign _T_19146 = _T_19145 | _T_19099; // @[Mux.scala 19:72:@15534.4]
  assign _T_19147 = _T_19146 | _T_19116; // @[Mux.scala 19:72:@15535.4]
  assign _T_19148 = _T_19147 | _T_19133; // @[Mux.scala 19:72:@15536.4]
  assign _T_19726 = {conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0}; // @[Mux.scala 19:72:@15886.4]
  assign _T_19733 = {conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8}; // @[Mux.scala 19:72:@15893.4]
  assign _T_19734 = {conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,_T_19726}; // @[Mux.scala 19:72:@15894.4]
  assign _T_19736 = _T_2697 ? _T_19734 : 16'h0; // @[Mux.scala 19:72:@15895.4]
  assign _T_19743 = {conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1}; // @[Mux.scala 19:72:@15902.4]
  assign _T_19750 = {conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9}; // @[Mux.scala 19:72:@15909.4]
  assign _T_19751 = {conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,_T_19743}; // @[Mux.scala 19:72:@15910.4]
  assign _T_19753 = _T_2698 ? _T_19751 : 16'h0; // @[Mux.scala 19:72:@15911.4]
  assign _T_19760 = {conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2}; // @[Mux.scala 19:72:@15918.4]
  assign _T_19767 = {conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10}; // @[Mux.scala 19:72:@15925.4]
  assign _T_19768 = {conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,_T_19760}; // @[Mux.scala 19:72:@15926.4]
  assign _T_19770 = _T_2699 ? _T_19768 : 16'h0; // @[Mux.scala 19:72:@15927.4]
  assign _T_19777 = {conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3}; // @[Mux.scala 19:72:@15934.4]
  assign _T_19784 = {conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11}; // @[Mux.scala 19:72:@15941.4]
  assign _T_19785 = {conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,_T_19777}; // @[Mux.scala 19:72:@15942.4]
  assign _T_19787 = _T_2700 ? _T_19785 : 16'h0; // @[Mux.scala 19:72:@15943.4]
  assign _T_19794 = {conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4}; // @[Mux.scala 19:72:@15950.4]
  assign _T_19801 = {conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12}; // @[Mux.scala 19:72:@15957.4]
  assign _T_19802 = {conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,_T_19794}; // @[Mux.scala 19:72:@15958.4]
  assign _T_19804 = _T_2701 ? _T_19802 : 16'h0; // @[Mux.scala 19:72:@15959.4]
  assign _T_19811 = {conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5}; // @[Mux.scala 19:72:@15966.4]
  assign _T_19818 = {conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13}; // @[Mux.scala 19:72:@15973.4]
  assign _T_19819 = {conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,_T_19811}; // @[Mux.scala 19:72:@15974.4]
  assign _T_19821 = _T_2702 ? _T_19819 : 16'h0; // @[Mux.scala 19:72:@15975.4]
  assign _T_19828 = {conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6}; // @[Mux.scala 19:72:@15982.4]
  assign _T_19835 = {conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14}; // @[Mux.scala 19:72:@15989.4]
  assign _T_19836 = {conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,_T_19828}; // @[Mux.scala 19:72:@15990.4]
  assign _T_19838 = _T_2703 ? _T_19836 : 16'h0; // @[Mux.scala 19:72:@15991.4]
  assign _T_19845 = {conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7}; // @[Mux.scala 19:72:@15998.4]
  assign _T_19852 = {conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15}; // @[Mux.scala 19:72:@16005.4]
  assign _T_19853 = {conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,_T_19845}; // @[Mux.scala 19:72:@16006.4]
  assign _T_19855 = _T_2704 ? _T_19853 : 16'h0; // @[Mux.scala 19:72:@16007.4]
  assign _T_19870 = {conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,_T_19733}; // @[Mux.scala 19:72:@16022.4]
  assign _T_19872 = _T_2705 ? _T_19870 : 16'h0; // @[Mux.scala 19:72:@16023.4]
  assign _T_19887 = {conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,_T_19750}; // @[Mux.scala 19:72:@16038.4]
  assign _T_19889 = _T_2706 ? _T_19887 : 16'h0; // @[Mux.scala 19:72:@16039.4]
  assign _T_19904 = {conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,_T_19767}; // @[Mux.scala 19:72:@16054.4]
  assign _T_19906 = _T_2707 ? _T_19904 : 16'h0; // @[Mux.scala 19:72:@16055.4]
  assign _T_19921 = {conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,_T_19784}; // @[Mux.scala 19:72:@16070.4]
  assign _T_19923 = _T_2708 ? _T_19921 : 16'h0; // @[Mux.scala 19:72:@16071.4]
  assign _T_19938 = {conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,_T_19801}; // @[Mux.scala 19:72:@16086.4]
  assign _T_19940 = _T_2709 ? _T_19938 : 16'h0; // @[Mux.scala 19:72:@16087.4]
  assign _T_19955 = {conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,_T_19818}; // @[Mux.scala 19:72:@16102.4]
  assign _T_19957 = _T_2710 ? _T_19955 : 16'h0; // @[Mux.scala 19:72:@16103.4]
  assign _T_19972 = {conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,_T_19835}; // @[Mux.scala 19:72:@16118.4]
  assign _T_19974 = _T_2711 ? _T_19972 : 16'h0; // @[Mux.scala 19:72:@16119.4]
  assign _T_19989 = {conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,_T_19852}; // @[Mux.scala 19:72:@16134.4]
  assign _T_19991 = _T_2712 ? _T_19989 : 16'h0; // @[Mux.scala 19:72:@16135.4]
  assign _T_19992 = _T_19736 | _T_19753; // @[Mux.scala 19:72:@16136.4]
  assign _T_19993 = _T_19992 | _T_19770; // @[Mux.scala 19:72:@16137.4]
  assign _T_19994 = _T_19993 | _T_19787; // @[Mux.scala 19:72:@16138.4]
  assign _T_19995 = _T_19994 | _T_19804; // @[Mux.scala 19:72:@16139.4]
  assign _T_19996 = _T_19995 | _T_19821; // @[Mux.scala 19:72:@16140.4]
  assign _T_19997 = _T_19996 | _T_19838; // @[Mux.scala 19:72:@16141.4]
  assign _T_19998 = _T_19997 | _T_19855; // @[Mux.scala 19:72:@16142.4]
  assign _T_19999 = _T_19998 | _T_19872; // @[Mux.scala 19:72:@16143.4]
  assign _T_20000 = _T_19999 | _T_19889; // @[Mux.scala 19:72:@16144.4]
  assign _T_20001 = _T_20000 | _T_19906; // @[Mux.scala 19:72:@16145.4]
  assign _T_20002 = _T_20001 | _T_19923; // @[Mux.scala 19:72:@16146.4]
  assign _T_20003 = _T_20002 | _T_19940; // @[Mux.scala 19:72:@16147.4]
  assign _T_20004 = _T_20003 | _T_19957; // @[Mux.scala 19:72:@16148.4]
  assign _T_20005 = _T_20004 | _T_19974; // @[Mux.scala 19:72:@16149.4]
  assign _T_20006 = _T_20005 | _T_19991; // @[Mux.scala 19:72:@16150.4]
  assign _T_20584 = {conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0}; // @[Mux.scala 19:72:@16500.4]
  assign _T_20591 = {conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8}; // @[Mux.scala 19:72:@16507.4]
  assign _T_20592 = {conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,_T_20584}; // @[Mux.scala 19:72:@16508.4]
  assign _T_20594 = _T_2697 ? _T_20592 : 16'h0; // @[Mux.scala 19:72:@16509.4]
  assign _T_20601 = {conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1}; // @[Mux.scala 19:72:@16516.4]
  assign _T_20608 = {conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9}; // @[Mux.scala 19:72:@16523.4]
  assign _T_20609 = {conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,_T_20601}; // @[Mux.scala 19:72:@16524.4]
  assign _T_20611 = _T_2698 ? _T_20609 : 16'h0; // @[Mux.scala 19:72:@16525.4]
  assign _T_20618 = {conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2}; // @[Mux.scala 19:72:@16532.4]
  assign _T_20625 = {conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10}; // @[Mux.scala 19:72:@16539.4]
  assign _T_20626 = {conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,_T_20618}; // @[Mux.scala 19:72:@16540.4]
  assign _T_20628 = _T_2699 ? _T_20626 : 16'h0; // @[Mux.scala 19:72:@16541.4]
  assign _T_20635 = {conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3}; // @[Mux.scala 19:72:@16548.4]
  assign _T_20642 = {conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11}; // @[Mux.scala 19:72:@16555.4]
  assign _T_20643 = {conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,_T_20635}; // @[Mux.scala 19:72:@16556.4]
  assign _T_20645 = _T_2700 ? _T_20643 : 16'h0; // @[Mux.scala 19:72:@16557.4]
  assign _T_20652 = {conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4}; // @[Mux.scala 19:72:@16564.4]
  assign _T_20659 = {conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12}; // @[Mux.scala 19:72:@16571.4]
  assign _T_20660 = {conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,_T_20652}; // @[Mux.scala 19:72:@16572.4]
  assign _T_20662 = _T_2701 ? _T_20660 : 16'h0; // @[Mux.scala 19:72:@16573.4]
  assign _T_20669 = {conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5}; // @[Mux.scala 19:72:@16580.4]
  assign _T_20676 = {conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13}; // @[Mux.scala 19:72:@16587.4]
  assign _T_20677 = {conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,_T_20669}; // @[Mux.scala 19:72:@16588.4]
  assign _T_20679 = _T_2702 ? _T_20677 : 16'h0; // @[Mux.scala 19:72:@16589.4]
  assign _T_20686 = {conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6}; // @[Mux.scala 19:72:@16596.4]
  assign _T_20693 = {conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14}; // @[Mux.scala 19:72:@16603.4]
  assign _T_20694 = {conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,_T_20686}; // @[Mux.scala 19:72:@16604.4]
  assign _T_20696 = _T_2703 ? _T_20694 : 16'h0; // @[Mux.scala 19:72:@16605.4]
  assign _T_20703 = {conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7}; // @[Mux.scala 19:72:@16612.4]
  assign _T_20710 = {conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15}; // @[Mux.scala 19:72:@16619.4]
  assign _T_20711 = {conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,_T_20703}; // @[Mux.scala 19:72:@16620.4]
  assign _T_20713 = _T_2704 ? _T_20711 : 16'h0; // @[Mux.scala 19:72:@16621.4]
  assign _T_20728 = {conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,_T_20591}; // @[Mux.scala 19:72:@16636.4]
  assign _T_20730 = _T_2705 ? _T_20728 : 16'h0; // @[Mux.scala 19:72:@16637.4]
  assign _T_20745 = {conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,_T_20608}; // @[Mux.scala 19:72:@16652.4]
  assign _T_20747 = _T_2706 ? _T_20745 : 16'h0; // @[Mux.scala 19:72:@16653.4]
  assign _T_20762 = {conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,_T_20625}; // @[Mux.scala 19:72:@16668.4]
  assign _T_20764 = _T_2707 ? _T_20762 : 16'h0; // @[Mux.scala 19:72:@16669.4]
  assign _T_20779 = {conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,_T_20642}; // @[Mux.scala 19:72:@16684.4]
  assign _T_20781 = _T_2708 ? _T_20779 : 16'h0; // @[Mux.scala 19:72:@16685.4]
  assign _T_20796 = {conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,_T_20659}; // @[Mux.scala 19:72:@16700.4]
  assign _T_20798 = _T_2709 ? _T_20796 : 16'h0; // @[Mux.scala 19:72:@16701.4]
  assign _T_20813 = {conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,_T_20676}; // @[Mux.scala 19:72:@16716.4]
  assign _T_20815 = _T_2710 ? _T_20813 : 16'h0; // @[Mux.scala 19:72:@16717.4]
  assign _T_20830 = {conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,_T_20693}; // @[Mux.scala 19:72:@16732.4]
  assign _T_20832 = _T_2711 ? _T_20830 : 16'h0; // @[Mux.scala 19:72:@16733.4]
  assign _T_20847 = {conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,_T_20710}; // @[Mux.scala 19:72:@16748.4]
  assign _T_20849 = _T_2712 ? _T_20847 : 16'h0; // @[Mux.scala 19:72:@16749.4]
  assign _T_20850 = _T_20594 | _T_20611; // @[Mux.scala 19:72:@16750.4]
  assign _T_20851 = _T_20850 | _T_20628; // @[Mux.scala 19:72:@16751.4]
  assign _T_20852 = _T_20851 | _T_20645; // @[Mux.scala 19:72:@16752.4]
  assign _T_20853 = _T_20852 | _T_20662; // @[Mux.scala 19:72:@16753.4]
  assign _T_20854 = _T_20853 | _T_20679; // @[Mux.scala 19:72:@16754.4]
  assign _T_20855 = _T_20854 | _T_20696; // @[Mux.scala 19:72:@16755.4]
  assign _T_20856 = _T_20855 | _T_20713; // @[Mux.scala 19:72:@16756.4]
  assign _T_20857 = _T_20856 | _T_20730; // @[Mux.scala 19:72:@16757.4]
  assign _T_20858 = _T_20857 | _T_20747; // @[Mux.scala 19:72:@16758.4]
  assign _T_20859 = _T_20858 | _T_20764; // @[Mux.scala 19:72:@16759.4]
  assign _T_20860 = _T_20859 | _T_20781; // @[Mux.scala 19:72:@16760.4]
  assign _T_20861 = _T_20860 | _T_20798; // @[Mux.scala 19:72:@16761.4]
  assign _T_20862 = _T_20861 | _T_20815; // @[Mux.scala 19:72:@16762.4]
  assign _T_20863 = _T_20862 | _T_20832; // @[Mux.scala 19:72:@16763.4]
  assign _T_20864 = _T_20863 | _T_20849; // @[Mux.scala 19:72:@16764.4]
  assign _T_21442 = {conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0}; // @[Mux.scala 19:72:@17114.4]
  assign _T_21449 = {conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8}; // @[Mux.scala 19:72:@17121.4]
  assign _T_21450 = {conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,_T_21442}; // @[Mux.scala 19:72:@17122.4]
  assign _T_21452 = _T_2697 ? _T_21450 : 16'h0; // @[Mux.scala 19:72:@17123.4]
  assign _T_21459 = {conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1}; // @[Mux.scala 19:72:@17130.4]
  assign _T_21466 = {conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9}; // @[Mux.scala 19:72:@17137.4]
  assign _T_21467 = {conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,_T_21459}; // @[Mux.scala 19:72:@17138.4]
  assign _T_21469 = _T_2698 ? _T_21467 : 16'h0; // @[Mux.scala 19:72:@17139.4]
  assign _T_21476 = {conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2}; // @[Mux.scala 19:72:@17146.4]
  assign _T_21483 = {conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10}; // @[Mux.scala 19:72:@17153.4]
  assign _T_21484 = {conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,_T_21476}; // @[Mux.scala 19:72:@17154.4]
  assign _T_21486 = _T_2699 ? _T_21484 : 16'h0; // @[Mux.scala 19:72:@17155.4]
  assign _T_21493 = {conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3}; // @[Mux.scala 19:72:@17162.4]
  assign _T_21500 = {conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11}; // @[Mux.scala 19:72:@17169.4]
  assign _T_21501 = {conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,_T_21493}; // @[Mux.scala 19:72:@17170.4]
  assign _T_21503 = _T_2700 ? _T_21501 : 16'h0; // @[Mux.scala 19:72:@17171.4]
  assign _T_21510 = {conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4}; // @[Mux.scala 19:72:@17178.4]
  assign _T_21517 = {conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12}; // @[Mux.scala 19:72:@17185.4]
  assign _T_21518 = {conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,_T_21510}; // @[Mux.scala 19:72:@17186.4]
  assign _T_21520 = _T_2701 ? _T_21518 : 16'h0; // @[Mux.scala 19:72:@17187.4]
  assign _T_21527 = {conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5}; // @[Mux.scala 19:72:@17194.4]
  assign _T_21534 = {conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13}; // @[Mux.scala 19:72:@17201.4]
  assign _T_21535 = {conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,_T_21527}; // @[Mux.scala 19:72:@17202.4]
  assign _T_21537 = _T_2702 ? _T_21535 : 16'h0; // @[Mux.scala 19:72:@17203.4]
  assign _T_21544 = {conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6}; // @[Mux.scala 19:72:@17210.4]
  assign _T_21551 = {conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14}; // @[Mux.scala 19:72:@17217.4]
  assign _T_21552 = {conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,_T_21544}; // @[Mux.scala 19:72:@17218.4]
  assign _T_21554 = _T_2703 ? _T_21552 : 16'h0; // @[Mux.scala 19:72:@17219.4]
  assign _T_21561 = {conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7}; // @[Mux.scala 19:72:@17226.4]
  assign _T_21568 = {conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15}; // @[Mux.scala 19:72:@17233.4]
  assign _T_21569 = {conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,_T_21561}; // @[Mux.scala 19:72:@17234.4]
  assign _T_21571 = _T_2704 ? _T_21569 : 16'h0; // @[Mux.scala 19:72:@17235.4]
  assign _T_21586 = {conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,_T_21449}; // @[Mux.scala 19:72:@17250.4]
  assign _T_21588 = _T_2705 ? _T_21586 : 16'h0; // @[Mux.scala 19:72:@17251.4]
  assign _T_21603 = {conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,_T_21466}; // @[Mux.scala 19:72:@17266.4]
  assign _T_21605 = _T_2706 ? _T_21603 : 16'h0; // @[Mux.scala 19:72:@17267.4]
  assign _T_21620 = {conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,_T_21483}; // @[Mux.scala 19:72:@17282.4]
  assign _T_21622 = _T_2707 ? _T_21620 : 16'h0; // @[Mux.scala 19:72:@17283.4]
  assign _T_21637 = {conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,_T_21500}; // @[Mux.scala 19:72:@17298.4]
  assign _T_21639 = _T_2708 ? _T_21637 : 16'h0; // @[Mux.scala 19:72:@17299.4]
  assign _T_21654 = {conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,_T_21517}; // @[Mux.scala 19:72:@17314.4]
  assign _T_21656 = _T_2709 ? _T_21654 : 16'h0; // @[Mux.scala 19:72:@17315.4]
  assign _T_21671 = {conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,_T_21534}; // @[Mux.scala 19:72:@17330.4]
  assign _T_21673 = _T_2710 ? _T_21671 : 16'h0; // @[Mux.scala 19:72:@17331.4]
  assign _T_21688 = {conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,_T_21551}; // @[Mux.scala 19:72:@17346.4]
  assign _T_21690 = _T_2711 ? _T_21688 : 16'h0; // @[Mux.scala 19:72:@17347.4]
  assign _T_21705 = {conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,_T_21568}; // @[Mux.scala 19:72:@17362.4]
  assign _T_21707 = _T_2712 ? _T_21705 : 16'h0; // @[Mux.scala 19:72:@17363.4]
  assign _T_21708 = _T_21452 | _T_21469; // @[Mux.scala 19:72:@17364.4]
  assign _T_21709 = _T_21708 | _T_21486; // @[Mux.scala 19:72:@17365.4]
  assign _T_21710 = _T_21709 | _T_21503; // @[Mux.scala 19:72:@17366.4]
  assign _T_21711 = _T_21710 | _T_21520; // @[Mux.scala 19:72:@17367.4]
  assign _T_21712 = _T_21711 | _T_21537; // @[Mux.scala 19:72:@17368.4]
  assign _T_21713 = _T_21712 | _T_21554; // @[Mux.scala 19:72:@17369.4]
  assign _T_21714 = _T_21713 | _T_21571; // @[Mux.scala 19:72:@17370.4]
  assign _T_21715 = _T_21714 | _T_21588; // @[Mux.scala 19:72:@17371.4]
  assign _T_21716 = _T_21715 | _T_21605; // @[Mux.scala 19:72:@17372.4]
  assign _T_21717 = _T_21716 | _T_21622; // @[Mux.scala 19:72:@17373.4]
  assign _T_21718 = _T_21717 | _T_21639; // @[Mux.scala 19:72:@17374.4]
  assign _T_21719 = _T_21718 | _T_21656; // @[Mux.scala 19:72:@17375.4]
  assign _T_21720 = _T_21719 | _T_21673; // @[Mux.scala 19:72:@17376.4]
  assign _T_21721 = _T_21720 | _T_21690; // @[Mux.scala 19:72:@17377.4]
  assign _T_21722 = _T_21721 | _T_21707; // @[Mux.scala 19:72:@17378.4]
  assign _T_22300 = {conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0}; // @[Mux.scala 19:72:@17728.4]
  assign _T_22307 = {conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8}; // @[Mux.scala 19:72:@17735.4]
  assign _T_22308 = {conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,_T_22300}; // @[Mux.scala 19:72:@17736.4]
  assign _T_22310 = _T_2697 ? _T_22308 : 16'h0; // @[Mux.scala 19:72:@17737.4]
  assign _T_22317 = {conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1}; // @[Mux.scala 19:72:@17744.4]
  assign _T_22324 = {conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9}; // @[Mux.scala 19:72:@17751.4]
  assign _T_22325 = {conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,_T_22317}; // @[Mux.scala 19:72:@17752.4]
  assign _T_22327 = _T_2698 ? _T_22325 : 16'h0; // @[Mux.scala 19:72:@17753.4]
  assign _T_22334 = {conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2}; // @[Mux.scala 19:72:@17760.4]
  assign _T_22341 = {conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10}; // @[Mux.scala 19:72:@17767.4]
  assign _T_22342 = {conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,_T_22334}; // @[Mux.scala 19:72:@17768.4]
  assign _T_22344 = _T_2699 ? _T_22342 : 16'h0; // @[Mux.scala 19:72:@17769.4]
  assign _T_22351 = {conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3}; // @[Mux.scala 19:72:@17776.4]
  assign _T_22358 = {conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11}; // @[Mux.scala 19:72:@17783.4]
  assign _T_22359 = {conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,_T_22351}; // @[Mux.scala 19:72:@17784.4]
  assign _T_22361 = _T_2700 ? _T_22359 : 16'h0; // @[Mux.scala 19:72:@17785.4]
  assign _T_22368 = {conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4}; // @[Mux.scala 19:72:@17792.4]
  assign _T_22375 = {conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12}; // @[Mux.scala 19:72:@17799.4]
  assign _T_22376 = {conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,_T_22368}; // @[Mux.scala 19:72:@17800.4]
  assign _T_22378 = _T_2701 ? _T_22376 : 16'h0; // @[Mux.scala 19:72:@17801.4]
  assign _T_22385 = {conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5}; // @[Mux.scala 19:72:@17808.4]
  assign _T_22392 = {conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13}; // @[Mux.scala 19:72:@17815.4]
  assign _T_22393 = {conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,_T_22385}; // @[Mux.scala 19:72:@17816.4]
  assign _T_22395 = _T_2702 ? _T_22393 : 16'h0; // @[Mux.scala 19:72:@17817.4]
  assign _T_22402 = {conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6}; // @[Mux.scala 19:72:@17824.4]
  assign _T_22409 = {conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14}; // @[Mux.scala 19:72:@17831.4]
  assign _T_22410 = {conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,_T_22402}; // @[Mux.scala 19:72:@17832.4]
  assign _T_22412 = _T_2703 ? _T_22410 : 16'h0; // @[Mux.scala 19:72:@17833.4]
  assign _T_22419 = {conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7}; // @[Mux.scala 19:72:@17840.4]
  assign _T_22426 = {conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15}; // @[Mux.scala 19:72:@17847.4]
  assign _T_22427 = {conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,_T_22419}; // @[Mux.scala 19:72:@17848.4]
  assign _T_22429 = _T_2704 ? _T_22427 : 16'h0; // @[Mux.scala 19:72:@17849.4]
  assign _T_22444 = {conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,_T_22307}; // @[Mux.scala 19:72:@17864.4]
  assign _T_22446 = _T_2705 ? _T_22444 : 16'h0; // @[Mux.scala 19:72:@17865.4]
  assign _T_22461 = {conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,_T_22324}; // @[Mux.scala 19:72:@17880.4]
  assign _T_22463 = _T_2706 ? _T_22461 : 16'h0; // @[Mux.scala 19:72:@17881.4]
  assign _T_22478 = {conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,_T_22341}; // @[Mux.scala 19:72:@17896.4]
  assign _T_22480 = _T_2707 ? _T_22478 : 16'h0; // @[Mux.scala 19:72:@17897.4]
  assign _T_22495 = {conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,_T_22358}; // @[Mux.scala 19:72:@17912.4]
  assign _T_22497 = _T_2708 ? _T_22495 : 16'h0; // @[Mux.scala 19:72:@17913.4]
  assign _T_22512 = {conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,_T_22375}; // @[Mux.scala 19:72:@17928.4]
  assign _T_22514 = _T_2709 ? _T_22512 : 16'h0; // @[Mux.scala 19:72:@17929.4]
  assign _T_22529 = {conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,_T_22392}; // @[Mux.scala 19:72:@17944.4]
  assign _T_22531 = _T_2710 ? _T_22529 : 16'h0; // @[Mux.scala 19:72:@17945.4]
  assign _T_22546 = {conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,_T_22409}; // @[Mux.scala 19:72:@17960.4]
  assign _T_22548 = _T_2711 ? _T_22546 : 16'h0; // @[Mux.scala 19:72:@17961.4]
  assign _T_22563 = {conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,_T_22426}; // @[Mux.scala 19:72:@17976.4]
  assign _T_22565 = _T_2712 ? _T_22563 : 16'h0; // @[Mux.scala 19:72:@17977.4]
  assign _T_22566 = _T_22310 | _T_22327; // @[Mux.scala 19:72:@17978.4]
  assign _T_22567 = _T_22566 | _T_22344; // @[Mux.scala 19:72:@17979.4]
  assign _T_22568 = _T_22567 | _T_22361; // @[Mux.scala 19:72:@17980.4]
  assign _T_22569 = _T_22568 | _T_22378; // @[Mux.scala 19:72:@17981.4]
  assign _T_22570 = _T_22569 | _T_22395; // @[Mux.scala 19:72:@17982.4]
  assign _T_22571 = _T_22570 | _T_22412; // @[Mux.scala 19:72:@17983.4]
  assign _T_22572 = _T_22571 | _T_22429; // @[Mux.scala 19:72:@17984.4]
  assign _T_22573 = _T_22572 | _T_22446; // @[Mux.scala 19:72:@17985.4]
  assign _T_22574 = _T_22573 | _T_22463; // @[Mux.scala 19:72:@17986.4]
  assign _T_22575 = _T_22574 | _T_22480; // @[Mux.scala 19:72:@17987.4]
  assign _T_22576 = _T_22575 | _T_22497; // @[Mux.scala 19:72:@17988.4]
  assign _T_22577 = _T_22576 | _T_22514; // @[Mux.scala 19:72:@17989.4]
  assign _T_22578 = _T_22577 | _T_22531; // @[Mux.scala 19:72:@17990.4]
  assign _T_22579 = _T_22578 | _T_22548; // @[Mux.scala 19:72:@17991.4]
  assign _T_22580 = _T_22579 | _T_22565; // @[Mux.scala 19:72:@17992.4]
  assign _T_23158 = {conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0}; // @[Mux.scala 19:72:@18342.4]
  assign _T_23165 = {conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8}; // @[Mux.scala 19:72:@18349.4]
  assign _T_23166 = {conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,_T_23158}; // @[Mux.scala 19:72:@18350.4]
  assign _T_23168 = _T_2697 ? _T_23166 : 16'h0; // @[Mux.scala 19:72:@18351.4]
  assign _T_23175 = {conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1}; // @[Mux.scala 19:72:@18358.4]
  assign _T_23182 = {conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9}; // @[Mux.scala 19:72:@18365.4]
  assign _T_23183 = {conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,_T_23175}; // @[Mux.scala 19:72:@18366.4]
  assign _T_23185 = _T_2698 ? _T_23183 : 16'h0; // @[Mux.scala 19:72:@18367.4]
  assign _T_23192 = {conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2}; // @[Mux.scala 19:72:@18374.4]
  assign _T_23199 = {conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10}; // @[Mux.scala 19:72:@18381.4]
  assign _T_23200 = {conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,_T_23192}; // @[Mux.scala 19:72:@18382.4]
  assign _T_23202 = _T_2699 ? _T_23200 : 16'h0; // @[Mux.scala 19:72:@18383.4]
  assign _T_23209 = {conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3}; // @[Mux.scala 19:72:@18390.4]
  assign _T_23216 = {conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11}; // @[Mux.scala 19:72:@18397.4]
  assign _T_23217 = {conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,_T_23209}; // @[Mux.scala 19:72:@18398.4]
  assign _T_23219 = _T_2700 ? _T_23217 : 16'h0; // @[Mux.scala 19:72:@18399.4]
  assign _T_23226 = {conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4}; // @[Mux.scala 19:72:@18406.4]
  assign _T_23233 = {conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12}; // @[Mux.scala 19:72:@18413.4]
  assign _T_23234 = {conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,_T_23226}; // @[Mux.scala 19:72:@18414.4]
  assign _T_23236 = _T_2701 ? _T_23234 : 16'h0; // @[Mux.scala 19:72:@18415.4]
  assign _T_23243 = {conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5}; // @[Mux.scala 19:72:@18422.4]
  assign _T_23250 = {conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13}; // @[Mux.scala 19:72:@18429.4]
  assign _T_23251 = {conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,_T_23243}; // @[Mux.scala 19:72:@18430.4]
  assign _T_23253 = _T_2702 ? _T_23251 : 16'h0; // @[Mux.scala 19:72:@18431.4]
  assign _T_23260 = {conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6}; // @[Mux.scala 19:72:@18438.4]
  assign _T_23267 = {conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14}; // @[Mux.scala 19:72:@18445.4]
  assign _T_23268 = {conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,_T_23260}; // @[Mux.scala 19:72:@18446.4]
  assign _T_23270 = _T_2703 ? _T_23268 : 16'h0; // @[Mux.scala 19:72:@18447.4]
  assign _T_23277 = {conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7}; // @[Mux.scala 19:72:@18454.4]
  assign _T_23284 = {conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15}; // @[Mux.scala 19:72:@18461.4]
  assign _T_23285 = {conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,_T_23277}; // @[Mux.scala 19:72:@18462.4]
  assign _T_23287 = _T_2704 ? _T_23285 : 16'h0; // @[Mux.scala 19:72:@18463.4]
  assign _T_23302 = {conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,_T_23165}; // @[Mux.scala 19:72:@18478.4]
  assign _T_23304 = _T_2705 ? _T_23302 : 16'h0; // @[Mux.scala 19:72:@18479.4]
  assign _T_23319 = {conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,_T_23182}; // @[Mux.scala 19:72:@18494.4]
  assign _T_23321 = _T_2706 ? _T_23319 : 16'h0; // @[Mux.scala 19:72:@18495.4]
  assign _T_23336 = {conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,_T_23199}; // @[Mux.scala 19:72:@18510.4]
  assign _T_23338 = _T_2707 ? _T_23336 : 16'h0; // @[Mux.scala 19:72:@18511.4]
  assign _T_23353 = {conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,_T_23216}; // @[Mux.scala 19:72:@18526.4]
  assign _T_23355 = _T_2708 ? _T_23353 : 16'h0; // @[Mux.scala 19:72:@18527.4]
  assign _T_23370 = {conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,_T_23233}; // @[Mux.scala 19:72:@18542.4]
  assign _T_23372 = _T_2709 ? _T_23370 : 16'h0; // @[Mux.scala 19:72:@18543.4]
  assign _T_23387 = {conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,_T_23250}; // @[Mux.scala 19:72:@18558.4]
  assign _T_23389 = _T_2710 ? _T_23387 : 16'h0; // @[Mux.scala 19:72:@18559.4]
  assign _T_23404 = {conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,_T_23267}; // @[Mux.scala 19:72:@18574.4]
  assign _T_23406 = _T_2711 ? _T_23404 : 16'h0; // @[Mux.scala 19:72:@18575.4]
  assign _T_23421 = {conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,_T_23284}; // @[Mux.scala 19:72:@18590.4]
  assign _T_23423 = _T_2712 ? _T_23421 : 16'h0; // @[Mux.scala 19:72:@18591.4]
  assign _T_23424 = _T_23168 | _T_23185; // @[Mux.scala 19:72:@18592.4]
  assign _T_23425 = _T_23424 | _T_23202; // @[Mux.scala 19:72:@18593.4]
  assign _T_23426 = _T_23425 | _T_23219; // @[Mux.scala 19:72:@18594.4]
  assign _T_23427 = _T_23426 | _T_23236; // @[Mux.scala 19:72:@18595.4]
  assign _T_23428 = _T_23427 | _T_23253; // @[Mux.scala 19:72:@18596.4]
  assign _T_23429 = _T_23428 | _T_23270; // @[Mux.scala 19:72:@18597.4]
  assign _T_23430 = _T_23429 | _T_23287; // @[Mux.scala 19:72:@18598.4]
  assign _T_23431 = _T_23430 | _T_23304; // @[Mux.scala 19:72:@18599.4]
  assign _T_23432 = _T_23431 | _T_23321; // @[Mux.scala 19:72:@18600.4]
  assign _T_23433 = _T_23432 | _T_23338; // @[Mux.scala 19:72:@18601.4]
  assign _T_23434 = _T_23433 | _T_23355; // @[Mux.scala 19:72:@18602.4]
  assign _T_23435 = _T_23434 | _T_23372; // @[Mux.scala 19:72:@18603.4]
  assign _T_23436 = _T_23435 | _T_23389; // @[Mux.scala 19:72:@18604.4]
  assign _T_23437 = _T_23436 | _T_23406; // @[Mux.scala 19:72:@18605.4]
  assign _T_23438 = _T_23437 | _T_23423; // @[Mux.scala 19:72:@18606.4]
  assign _T_24016 = {conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0}; // @[Mux.scala 19:72:@18956.4]
  assign _T_24023 = {conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8}; // @[Mux.scala 19:72:@18963.4]
  assign _T_24024 = {conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,_T_24016}; // @[Mux.scala 19:72:@18964.4]
  assign _T_24026 = _T_2697 ? _T_24024 : 16'h0; // @[Mux.scala 19:72:@18965.4]
  assign _T_24033 = {conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1}; // @[Mux.scala 19:72:@18972.4]
  assign _T_24040 = {conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9}; // @[Mux.scala 19:72:@18979.4]
  assign _T_24041 = {conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,_T_24033}; // @[Mux.scala 19:72:@18980.4]
  assign _T_24043 = _T_2698 ? _T_24041 : 16'h0; // @[Mux.scala 19:72:@18981.4]
  assign _T_24050 = {conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2}; // @[Mux.scala 19:72:@18988.4]
  assign _T_24057 = {conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10}; // @[Mux.scala 19:72:@18995.4]
  assign _T_24058 = {conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,_T_24050}; // @[Mux.scala 19:72:@18996.4]
  assign _T_24060 = _T_2699 ? _T_24058 : 16'h0; // @[Mux.scala 19:72:@18997.4]
  assign _T_24067 = {conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3}; // @[Mux.scala 19:72:@19004.4]
  assign _T_24074 = {conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11}; // @[Mux.scala 19:72:@19011.4]
  assign _T_24075 = {conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,_T_24067}; // @[Mux.scala 19:72:@19012.4]
  assign _T_24077 = _T_2700 ? _T_24075 : 16'h0; // @[Mux.scala 19:72:@19013.4]
  assign _T_24084 = {conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4}; // @[Mux.scala 19:72:@19020.4]
  assign _T_24091 = {conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12}; // @[Mux.scala 19:72:@19027.4]
  assign _T_24092 = {conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,_T_24084}; // @[Mux.scala 19:72:@19028.4]
  assign _T_24094 = _T_2701 ? _T_24092 : 16'h0; // @[Mux.scala 19:72:@19029.4]
  assign _T_24101 = {conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5}; // @[Mux.scala 19:72:@19036.4]
  assign _T_24108 = {conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13}; // @[Mux.scala 19:72:@19043.4]
  assign _T_24109 = {conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,_T_24101}; // @[Mux.scala 19:72:@19044.4]
  assign _T_24111 = _T_2702 ? _T_24109 : 16'h0; // @[Mux.scala 19:72:@19045.4]
  assign _T_24118 = {conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6}; // @[Mux.scala 19:72:@19052.4]
  assign _T_24125 = {conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14}; // @[Mux.scala 19:72:@19059.4]
  assign _T_24126 = {conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,_T_24118}; // @[Mux.scala 19:72:@19060.4]
  assign _T_24128 = _T_2703 ? _T_24126 : 16'h0; // @[Mux.scala 19:72:@19061.4]
  assign _T_24135 = {conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7}; // @[Mux.scala 19:72:@19068.4]
  assign _T_24142 = {conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15}; // @[Mux.scala 19:72:@19075.4]
  assign _T_24143 = {conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,_T_24135}; // @[Mux.scala 19:72:@19076.4]
  assign _T_24145 = _T_2704 ? _T_24143 : 16'h0; // @[Mux.scala 19:72:@19077.4]
  assign _T_24160 = {conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,_T_24023}; // @[Mux.scala 19:72:@19092.4]
  assign _T_24162 = _T_2705 ? _T_24160 : 16'h0; // @[Mux.scala 19:72:@19093.4]
  assign _T_24177 = {conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,_T_24040}; // @[Mux.scala 19:72:@19108.4]
  assign _T_24179 = _T_2706 ? _T_24177 : 16'h0; // @[Mux.scala 19:72:@19109.4]
  assign _T_24194 = {conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,_T_24057}; // @[Mux.scala 19:72:@19124.4]
  assign _T_24196 = _T_2707 ? _T_24194 : 16'h0; // @[Mux.scala 19:72:@19125.4]
  assign _T_24211 = {conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,_T_24074}; // @[Mux.scala 19:72:@19140.4]
  assign _T_24213 = _T_2708 ? _T_24211 : 16'h0; // @[Mux.scala 19:72:@19141.4]
  assign _T_24228 = {conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,_T_24091}; // @[Mux.scala 19:72:@19156.4]
  assign _T_24230 = _T_2709 ? _T_24228 : 16'h0; // @[Mux.scala 19:72:@19157.4]
  assign _T_24245 = {conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,_T_24108}; // @[Mux.scala 19:72:@19172.4]
  assign _T_24247 = _T_2710 ? _T_24245 : 16'h0; // @[Mux.scala 19:72:@19173.4]
  assign _T_24262 = {conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,_T_24125}; // @[Mux.scala 19:72:@19188.4]
  assign _T_24264 = _T_2711 ? _T_24262 : 16'h0; // @[Mux.scala 19:72:@19189.4]
  assign _T_24279 = {conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,_T_24142}; // @[Mux.scala 19:72:@19204.4]
  assign _T_24281 = _T_2712 ? _T_24279 : 16'h0; // @[Mux.scala 19:72:@19205.4]
  assign _T_24282 = _T_24026 | _T_24043; // @[Mux.scala 19:72:@19206.4]
  assign _T_24283 = _T_24282 | _T_24060; // @[Mux.scala 19:72:@19207.4]
  assign _T_24284 = _T_24283 | _T_24077; // @[Mux.scala 19:72:@19208.4]
  assign _T_24285 = _T_24284 | _T_24094; // @[Mux.scala 19:72:@19209.4]
  assign _T_24286 = _T_24285 | _T_24111; // @[Mux.scala 19:72:@19210.4]
  assign _T_24287 = _T_24286 | _T_24128; // @[Mux.scala 19:72:@19211.4]
  assign _T_24288 = _T_24287 | _T_24145; // @[Mux.scala 19:72:@19212.4]
  assign _T_24289 = _T_24288 | _T_24162; // @[Mux.scala 19:72:@19213.4]
  assign _T_24290 = _T_24289 | _T_24179; // @[Mux.scala 19:72:@19214.4]
  assign _T_24291 = _T_24290 | _T_24196; // @[Mux.scala 19:72:@19215.4]
  assign _T_24292 = _T_24291 | _T_24213; // @[Mux.scala 19:72:@19216.4]
  assign _T_24293 = _T_24292 | _T_24230; // @[Mux.scala 19:72:@19217.4]
  assign _T_24294 = _T_24293 | _T_24247; // @[Mux.scala 19:72:@19218.4]
  assign _T_24295 = _T_24294 | _T_24264; // @[Mux.scala 19:72:@19219.4]
  assign _T_24296 = _T_24295 | _T_24281; // @[Mux.scala 19:72:@19220.4]
  assign _T_24874 = {conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0}; // @[Mux.scala 19:72:@19570.4]
  assign _T_24881 = {conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8}; // @[Mux.scala 19:72:@19577.4]
  assign _T_24882 = {conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,_T_24874}; // @[Mux.scala 19:72:@19578.4]
  assign _T_24884 = _T_2697 ? _T_24882 : 16'h0; // @[Mux.scala 19:72:@19579.4]
  assign _T_24891 = {conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1}; // @[Mux.scala 19:72:@19586.4]
  assign _T_24898 = {conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9}; // @[Mux.scala 19:72:@19593.4]
  assign _T_24899 = {conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,_T_24891}; // @[Mux.scala 19:72:@19594.4]
  assign _T_24901 = _T_2698 ? _T_24899 : 16'h0; // @[Mux.scala 19:72:@19595.4]
  assign _T_24908 = {conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2}; // @[Mux.scala 19:72:@19602.4]
  assign _T_24915 = {conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10}; // @[Mux.scala 19:72:@19609.4]
  assign _T_24916 = {conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,_T_24908}; // @[Mux.scala 19:72:@19610.4]
  assign _T_24918 = _T_2699 ? _T_24916 : 16'h0; // @[Mux.scala 19:72:@19611.4]
  assign _T_24925 = {conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3}; // @[Mux.scala 19:72:@19618.4]
  assign _T_24932 = {conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11}; // @[Mux.scala 19:72:@19625.4]
  assign _T_24933 = {conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,_T_24925}; // @[Mux.scala 19:72:@19626.4]
  assign _T_24935 = _T_2700 ? _T_24933 : 16'h0; // @[Mux.scala 19:72:@19627.4]
  assign _T_24942 = {conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4}; // @[Mux.scala 19:72:@19634.4]
  assign _T_24949 = {conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12}; // @[Mux.scala 19:72:@19641.4]
  assign _T_24950 = {conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,_T_24942}; // @[Mux.scala 19:72:@19642.4]
  assign _T_24952 = _T_2701 ? _T_24950 : 16'h0; // @[Mux.scala 19:72:@19643.4]
  assign _T_24959 = {conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5}; // @[Mux.scala 19:72:@19650.4]
  assign _T_24966 = {conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13}; // @[Mux.scala 19:72:@19657.4]
  assign _T_24967 = {conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,_T_24959}; // @[Mux.scala 19:72:@19658.4]
  assign _T_24969 = _T_2702 ? _T_24967 : 16'h0; // @[Mux.scala 19:72:@19659.4]
  assign _T_24976 = {conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6}; // @[Mux.scala 19:72:@19666.4]
  assign _T_24983 = {conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14}; // @[Mux.scala 19:72:@19673.4]
  assign _T_24984 = {conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,_T_24976}; // @[Mux.scala 19:72:@19674.4]
  assign _T_24986 = _T_2703 ? _T_24984 : 16'h0; // @[Mux.scala 19:72:@19675.4]
  assign _T_24993 = {conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7}; // @[Mux.scala 19:72:@19682.4]
  assign _T_25000 = {conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15}; // @[Mux.scala 19:72:@19689.4]
  assign _T_25001 = {conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,_T_24993}; // @[Mux.scala 19:72:@19690.4]
  assign _T_25003 = _T_2704 ? _T_25001 : 16'h0; // @[Mux.scala 19:72:@19691.4]
  assign _T_25018 = {conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,_T_24881}; // @[Mux.scala 19:72:@19706.4]
  assign _T_25020 = _T_2705 ? _T_25018 : 16'h0; // @[Mux.scala 19:72:@19707.4]
  assign _T_25035 = {conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,_T_24898}; // @[Mux.scala 19:72:@19722.4]
  assign _T_25037 = _T_2706 ? _T_25035 : 16'h0; // @[Mux.scala 19:72:@19723.4]
  assign _T_25052 = {conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,_T_24915}; // @[Mux.scala 19:72:@19738.4]
  assign _T_25054 = _T_2707 ? _T_25052 : 16'h0; // @[Mux.scala 19:72:@19739.4]
  assign _T_25069 = {conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,_T_24932}; // @[Mux.scala 19:72:@19754.4]
  assign _T_25071 = _T_2708 ? _T_25069 : 16'h0; // @[Mux.scala 19:72:@19755.4]
  assign _T_25086 = {conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,_T_24949}; // @[Mux.scala 19:72:@19770.4]
  assign _T_25088 = _T_2709 ? _T_25086 : 16'h0; // @[Mux.scala 19:72:@19771.4]
  assign _T_25103 = {conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,_T_24966}; // @[Mux.scala 19:72:@19786.4]
  assign _T_25105 = _T_2710 ? _T_25103 : 16'h0; // @[Mux.scala 19:72:@19787.4]
  assign _T_25120 = {conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,_T_24983}; // @[Mux.scala 19:72:@19802.4]
  assign _T_25122 = _T_2711 ? _T_25120 : 16'h0; // @[Mux.scala 19:72:@19803.4]
  assign _T_25137 = {conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,_T_25000}; // @[Mux.scala 19:72:@19818.4]
  assign _T_25139 = _T_2712 ? _T_25137 : 16'h0; // @[Mux.scala 19:72:@19819.4]
  assign _T_25140 = _T_24884 | _T_24901; // @[Mux.scala 19:72:@19820.4]
  assign _T_25141 = _T_25140 | _T_24918; // @[Mux.scala 19:72:@19821.4]
  assign _T_25142 = _T_25141 | _T_24935; // @[Mux.scala 19:72:@19822.4]
  assign _T_25143 = _T_25142 | _T_24952; // @[Mux.scala 19:72:@19823.4]
  assign _T_25144 = _T_25143 | _T_24969; // @[Mux.scala 19:72:@19824.4]
  assign _T_25145 = _T_25144 | _T_24986; // @[Mux.scala 19:72:@19825.4]
  assign _T_25146 = _T_25145 | _T_25003; // @[Mux.scala 19:72:@19826.4]
  assign _T_25147 = _T_25146 | _T_25020; // @[Mux.scala 19:72:@19827.4]
  assign _T_25148 = _T_25147 | _T_25037; // @[Mux.scala 19:72:@19828.4]
  assign _T_25149 = _T_25148 | _T_25054; // @[Mux.scala 19:72:@19829.4]
  assign _T_25150 = _T_25149 | _T_25071; // @[Mux.scala 19:72:@19830.4]
  assign _T_25151 = _T_25150 | _T_25088; // @[Mux.scala 19:72:@19831.4]
  assign _T_25152 = _T_25151 | _T_25105; // @[Mux.scala 19:72:@19832.4]
  assign _T_25153 = _T_25152 | _T_25122; // @[Mux.scala 19:72:@19833.4]
  assign _T_25154 = _T_25153 | _T_25139; // @[Mux.scala 19:72:@19834.4]
  assign _T_25732 = {conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0}; // @[Mux.scala 19:72:@20184.4]
  assign _T_25739 = {conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8}; // @[Mux.scala 19:72:@20191.4]
  assign _T_25740 = {conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,_T_25732}; // @[Mux.scala 19:72:@20192.4]
  assign _T_25742 = _T_2697 ? _T_25740 : 16'h0; // @[Mux.scala 19:72:@20193.4]
  assign _T_25749 = {conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1}; // @[Mux.scala 19:72:@20200.4]
  assign _T_25756 = {conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9}; // @[Mux.scala 19:72:@20207.4]
  assign _T_25757 = {conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,_T_25749}; // @[Mux.scala 19:72:@20208.4]
  assign _T_25759 = _T_2698 ? _T_25757 : 16'h0; // @[Mux.scala 19:72:@20209.4]
  assign _T_25766 = {conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2}; // @[Mux.scala 19:72:@20216.4]
  assign _T_25773 = {conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10}; // @[Mux.scala 19:72:@20223.4]
  assign _T_25774 = {conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,_T_25766}; // @[Mux.scala 19:72:@20224.4]
  assign _T_25776 = _T_2699 ? _T_25774 : 16'h0; // @[Mux.scala 19:72:@20225.4]
  assign _T_25783 = {conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3}; // @[Mux.scala 19:72:@20232.4]
  assign _T_25790 = {conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11}; // @[Mux.scala 19:72:@20239.4]
  assign _T_25791 = {conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,_T_25783}; // @[Mux.scala 19:72:@20240.4]
  assign _T_25793 = _T_2700 ? _T_25791 : 16'h0; // @[Mux.scala 19:72:@20241.4]
  assign _T_25800 = {conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4}; // @[Mux.scala 19:72:@20248.4]
  assign _T_25807 = {conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12}; // @[Mux.scala 19:72:@20255.4]
  assign _T_25808 = {conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,_T_25800}; // @[Mux.scala 19:72:@20256.4]
  assign _T_25810 = _T_2701 ? _T_25808 : 16'h0; // @[Mux.scala 19:72:@20257.4]
  assign _T_25817 = {conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5}; // @[Mux.scala 19:72:@20264.4]
  assign _T_25824 = {conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13}; // @[Mux.scala 19:72:@20271.4]
  assign _T_25825 = {conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,_T_25817}; // @[Mux.scala 19:72:@20272.4]
  assign _T_25827 = _T_2702 ? _T_25825 : 16'h0; // @[Mux.scala 19:72:@20273.4]
  assign _T_25834 = {conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6}; // @[Mux.scala 19:72:@20280.4]
  assign _T_25841 = {conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14}; // @[Mux.scala 19:72:@20287.4]
  assign _T_25842 = {conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,_T_25834}; // @[Mux.scala 19:72:@20288.4]
  assign _T_25844 = _T_2703 ? _T_25842 : 16'h0; // @[Mux.scala 19:72:@20289.4]
  assign _T_25851 = {conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7}; // @[Mux.scala 19:72:@20296.4]
  assign _T_25858 = {conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15}; // @[Mux.scala 19:72:@20303.4]
  assign _T_25859 = {conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,_T_25851}; // @[Mux.scala 19:72:@20304.4]
  assign _T_25861 = _T_2704 ? _T_25859 : 16'h0; // @[Mux.scala 19:72:@20305.4]
  assign _T_25876 = {conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,_T_25739}; // @[Mux.scala 19:72:@20320.4]
  assign _T_25878 = _T_2705 ? _T_25876 : 16'h0; // @[Mux.scala 19:72:@20321.4]
  assign _T_25893 = {conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,_T_25756}; // @[Mux.scala 19:72:@20336.4]
  assign _T_25895 = _T_2706 ? _T_25893 : 16'h0; // @[Mux.scala 19:72:@20337.4]
  assign _T_25910 = {conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,_T_25773}; // @[Mux.scala 19:72:@20352.4]
  assign _T_25912 = _T_2707 ? _T_25910 : 16'h0; // @[Mux.scala 19:72:@20353.4]
  assign _T_25927 = {conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,_T_25790}; // @[Mux.scala 19:72:@20368.4]
  assign _T_25929 = _T_2708 ? _T_25927 : 16'h0; // @[Mux.scala 19:72:@20369.4]
  assign _T_25944 = {conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,_T_25807}; // @[Mux.scala 19:72:@20384.4]
  assign _T_25946 = _T_2709 ? _T_25944 : 16'h0; // @[Mux.scala 19:72:@20385.4]
  assign _T_25961 = {conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,_T_25824}; // @[Mux.scala 19:72:@20400.4]
  assign _T_25963 = _T_2710 ? _T_25961 : 16'h0; // @[Mux.scala 19:72:@20401.4]
  assign _T_25978 = {conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,_T_25841}; // @[Mux.scala 19:72:@20416.4]
  assign _T_25980 = _T_2711 ? _T_25978 : 16'h0; // @[Mux.scala 19:72:@20417.4]
  assign _T_25995 = {conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,_T_25858}; // @[Mux.scala 19:72:@20432.4]
  assign _T_25997 = _T_2712 ? _T_25995 : 16'h0; // @[Mux.scala 19:72:@20433.4]
  assign _T_25998 = _T_25742 | _T_25759; // @[Mux.scala 19:72:@20434.4]
  assign _T_25999 = _T_25998 | _T_25776; // @[Mux.scala 19:72:@20435.4]
  assign _T_26000 = _T_25999 | _T_25793; // @[Mux.scala 19:72:@20436.4]
  assign _T_26001 = _T_26000 | _T_25810; // @[Mux.scala 19:72:@20437.4]
  assign _T_26002 = _T_26001 | _T_25827; // @[Mux.scala 19:72:@20438.4]
  assign _T_26003 = _T_26002 | _T_25844; // @[Mux.scala 19:72:@20439.4]
  assign _T_26004 = _T_26003 | _T_25861; // @[Mux.scala 19:72:@20440.4]
  assign _T_26005 = _T_26004 | _T_25878; // @[Mux.scala 19:72:@20441.4]
  assign _T_26006 = _T_26005 | _T_25895; // @[Mux.scala 19:72:@20442.4]
  assign _T_26007 = _T_26006 | _T_25912; // @[Mux.scala 19:72:@20443.4]
  assign _T_26008 = _T_26007 | _T_25929; // @[Mux.scala 19:72:@20444.4]
  assign _T_26009 = _T_26008 | _T_25946; // @[Mux.scala 19:72:@20445.4]
  assign _T_26010 = _T_26009 | _T_25963; // @[Mux.scala 19:72:@20446.4]
  assign _T_26011 = _T_26010 | _T_25980; // @[Mux.scala 19:72:@20447.4]
  assign _T_26012 = _T_26011 | _T_25997; // @[Mux.scala 19:72:@20448.4]
  assign _T_26590 = {conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0}; // @[Mux.scala 19:72:@20798.4]
  assign _T_26597 = {conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8}; // @[Mux.scala 19:72:@20805.4]
  assign _T_26598 = {conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,_T_26590}; // @[Mux.scala 19:72:@20806.4]
  assign _T_26600 = _T_2697 ? _T_26598 : 16'h0; // @[Mux.scala 19:72:@20807.4]
  assign _T_26607 = {conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1}; // @[Mux.scala 19:72:@20814.4]
  assign _T_26614 = {conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9}; // @[Mux.scala 19:72:@20821.4]
  assign _T_26615 = {conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,_T_26607}; // @[Mux.scala 19:72:@20822.4]
  assign _T_26617 = _T_2698 ? _T_26615 : 16'h0; // @[Mux.scala 19:72:@20823.4]
  assign _T_26624 = {conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2}; // @[Mux.scala 19:72:@20830.4]
  assign _T_26631 = {conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10}; // @[Mux.scala 19:72:@20837.4]
  assign _T_26632 = {conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,_T_26624}; // @[Mux.scala 19:72:@20838.4]
  assign _T_26634 = _T_2699 ? _T_26632 : 16'h0; // @[Mux.scala 19:72:@20839.4]
  assign _T_26641 = {conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3}; // @[Mux.scala 19:72:@20846.4]
  assign _T_26648 = {conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11}; // @[Mux.scala 19:72:@20853.4]
  assign _T_26649 = {conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,_T_26641}; // @[Mux.scala 19:72:@20854.4]
  assign _T_26651 = _T_2700 ? _T_26649 : 16'h0; // @[Mux.scala 19:72:@20855.4]
  assign _T_26658 = {conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4}; // @[Mux.scala 19:72:@20862.4]
  assign _T_26665 = {conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12}; // @[Mux.scala 19:72:@20869.4]
  assign _T_26666 = {conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,_T_26658}; // @[Mux.scala 19:72:@20870.4]
  assign _T_26668 = _T_2701 ? _T_26666 : 16'h0; // @[Mux.scala 19:72:@20871.4]
  assign _T_26675 = {conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5}; // @[Mux.scala 19:72:@20878.4]
  assign _T_26682 = {conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13}; // @[Mux.scala 19:72:@20885.4]
  assign _T_26683 = {conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,_T_26675}; // @[Mux.scala 19:72:@20886.4]
  assign _T_26685 = _T_2702 ? _T_26683 : 16'h0; // @[Mux.scala 19:72:@20887.4]
  assign _T_26692 = {conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6}; // @[Mux.scala 19:72:@20894.4]
  assign _T_26699 = {conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14}; // @[Mux.scala 19:72:@20901.4]
  assign _T_26700 = {conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,_T_26692}; // @[Mux.scala 19:72:@20902.4]
  assign _T_26702 = _T_2703 ? _T_26700 : 16'h0; // @[Mux.scala 19:72:@20903.4]
  assign _T_26709 = {conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7}; // @[Mux.scala 19:72:@20910.4]
  assign _T_26716 = {conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15}; // @[Mux.scala 19:72:@20917.4]
  assign _T_26717 = {conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,_T_26709}; // @[Mux.scala 19:72:@20918.4]
  assign _T_26719 = _T_2704 ? _T_26717 : 16'h0; // @[Mux.scala 19:72:@20919.4]
  assign _T_26734 = {conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,_T_26597}; // @[Mux.scala 19:72:@20934.4]
  assign _T_26736 = _T_2705 ? _T_26734 : 16'h0; // @[Mux.scala 19:72:@20935.4]
  assign _T_26751 = {conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,_T_26614}; // @[Mux.scala 19:72:@20950.4]
  assign _T_26753 = _T_2706 ? _T_26751 : 16'h0; // @[Mux.scala 19:72:@20951.4]
  assign _T_26768 = {conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,_T_26631}; // @[Mux.scala 19:72:@20966.4]
  assign _T_26770 = _T_2707 ? _T_26768 : 16'h0; // @[Mux.scala 19:72:@20967.4]
  assign _T_26785 = {conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,_T_26648}; // @[Mux.scala 19:72:@20982.4]
  assign _T_26787 = _T_2708 ? _T_26785 : 16'h0; // @[Mux.scala 19:72:@20983.4]
  assign _T_26802 = {conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,_T_26665}; // @[Mux.scala 19:72:@20998.4]
  assign _T_26804 = _T_2709 ? _T_26802 : 16'h0; // @[Mux.scala 19:72:@20999.4]
  assign _T_26819 = {conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,_T_26682}; // @[Mux.scala 19:72:@21014.4]
  assign _T_26821 = _T_2710 ? _T_26819 : 16'h0; // @[Mux.scala 19:72:@21015.4]
  assign _T_26836 = {conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,_T_26699}; // @[Mux.scala 19:72:@21030.4]
  assign _T_26838 = _T_2711 ? _T_26836 : 16'h0; // @[Mux.scala 19:72:@21031.4]
  assign _T_26853 = {conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,_T_26716}; // @[Mux.scala 19:72:@21046.4]
  assign _T_26855 = _T_2712 ? _T_26853 : 16'h0; // @[Mux.scala 19:72:@21047.4]
  assign _T_26856 = _T_26600 | _T_26617; // @[Mux.scala 19:72:@21048.4]
  assign _T_26857 = _T_26856 | _T_26634; // @[Mux.scala 19:72:@21049.4]
  assign _T_26858 = _T_26857 | _T_26651; // @[Mux.scala 19:72:@21050.4]
  assign _T_26859 = _T_26858 | _T_26668; // @[Mux.scala 19:72:@21051.4]
  assign _T_26860 = _T_26859 | _T_26685; // @[Mux.scala 19:72:@21052.4]
  assign _T_26861 = _T_26860 | _T_26702; // @[Mux.scala 19:72:@21053.4]
  assign _T_26862 = _T_26861 | _T_26719; // @[Mux.scala 19:72:@21054.4]
  assign _T_26863 = _T_26862 | _T_26736; // @[Mux.scala 19:72:@21055.4]
  assign _T_26864 = _T_26863 | _T_26753; // @[Mux.scala 19:72:@21056.4]
  assign _T_26865 = _T_26864 | _T_26770; // @[Mux.scala 19:72:@21057.4]
  assign _T_26866 = _T_26865 | _T_26787; // @[Mux.scala 19:72:@21058.4]
  assign _T_26867 = _T_26866 | _T_26804; // @[Mux.scala 19:72:@21059.4]
  assign _T_26868 = _T_26867 | _T_26821; // @[Mux.scala 19:72:@21060.4]
  assign _T_26869 = _T_26868 | _T_26838; // @[Mux.scala 19:72:@21061.4]
  assign _T_26870 = _T_26869 | _T_26855; // @[Mux.scala 19:72:@21062.4]
  assign _T_27448 = {conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0}; // @[Mux.scala 19:72:@21412.4]
  assign _T_27455 = {conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8}; // @[Mux.scala 19:72:@21419.4]
  assign _T_27456 = {conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,_T_27448}; // @[Mux.scala 19:72:@21420.4]
  assign _T_27458 = _T_2697 ? _T_27456 : 16'h0; // @[Mux.scala 19:72:@21421.4]
  assign _T_27465 = {conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1}; // @[Mux.scala 19:72:@21428.4]
  assign _T_27472 = {conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9}; // @[Mux.scala 19:72:@21435.4]
  assign _T_27473 = {conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,_T_27465}; // @[Mux.scala 19:72:@21436.4]
  assign _T_27475 = _T_2698 ? _T_27473 : 16'h0; // @[Mux.scala 19:72:@21437.4]
  assign _T_27482 = {conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2}; // @[Mux.scala 19:72:@21444.4]
  assign _T_27489 = {conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10}; // @[Mux.scala 19:72:@21451.4]
  assign _T_27490 = {conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,_T_27482}; // @[Mux.scala 19:72:@21452.4]
  assign _T_27492 = _T_2699 ? _T_27490 : 16'h0; // @[Mux.scala 19:72:@21453.4]
  assign _T_27499 = {conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3}; // @[Mux.scala 19:72:@21460.4]
  assign _T_27506 = {conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11}; // @[Mux.scala 19:72:@21467.4]
  assign _T_27507 = {conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,_T_27499}; // @[Mux.scala 19:72:@21468.4]
  assign _T_27509 = _T_2700 ? _T_27507 : 16'h0; // @[Mux.scala 19:72:@21469.4]
  assign _T_27516 = {conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4}; // @[Mux.scala 19:72:@21476.4]
  assign _T_27523 = {conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12}; // @[Mux.scala 19:72:@21483.4]
  assign _T_27524 = {conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,_T_27516}; // @[Mux.scala 19:72:@21484.4]
  assign _T_27526 = _T_2701 ? _T_27524 : 16'h0; // @[Mux.scala 19:72:@21485.4]
  assign _T_27533 = {conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5}; // @[Mux.scala 19:72:@21492.4]
  assign _T_27540 = {conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13}; // @[Mux.scala 19:72:@21499.4]
  assign _T_27541 = {conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,_T_27533}; // @[Mux.scala 19:72:@21500.4]
  assign _T_27543 = _T_2702 ? _T_27541 : 16'h0; // @[Mux.scala 19:72:@21501.4]
  assign _T_27550 = {conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6}; // @[Mux.scala 19:72:@21508.4]
  assign _T_27557 = {conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14}; // @[Mux.scala 19:72:@21515.4]
  assign _T_27558 = {conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,_T_27550}; // @[Mux.scala 19:72:@21516.4]
  assign _T_27560 = _T_2703 ? _T_27558 : 16'h0; // @[Mux.scala 19:72:@21517.4]
  assign _T_27567 = {conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7}; // @[Mux.scala 19:72:@21524.4]
  assign _T_27574 = {conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15}; // @[Mux.scala 19:72:@21531.4]
  assign _T_27575 = {conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,_T_27567}; // @[Mux.scala 19:72:@21532.4]
  assign _T_27577 = _T_2704 ? _T_27575 : 16'h0; // @[Mux.scala 19:72:@21533.4]
  assign _T_27592 = {conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,_T_27455}; // @[Mux.scala 19:72:@21548.4]
  assign _T_27594 = _T_2705 ? _T_27592 : 16'h0; // @[Mux.scala 19:72:@21549.4]
  assign _T_27609 = {conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,_T_27472}; // @[Mux.scala 19:72:@21564.4]
  assign _T_27611 = _T_2706 ? _T_27609 : 16'h0; // @[Mux.scala 19:72:@21565.4]
  assign _T_27626 = {conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,_T_27489}; // @[Mux.scala 19:72:@21580.4]
  assign _T_27628 = _T_2707 ? _T_27626 : 16'h0; // @[Mux.scala 19:72:@21581.4]
  assign _T_27643 = {conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,_T_27506}; // @[Mux.scala 19:72:@21596.4]
  assign _T_27645 = _T_2708 ? _T_27643 : 16'h0; // @[Mux.scala 19:72:@21597.4]
  assign _T_27660 = {conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,_T_27523}; // @[Mux.scala 19:72:@21612.4]
  assign _T_27662 = _T_2709 ? _T_27660 : 16'h0; // @[Mux.scala 19:72:@21613.4]
  assign _T_27677 = {conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,_T_27540}; // @[Mux.scala 19:72:@21628.4]
  assign _T_27679 = _T_2710 ? _T_27677 : 16'h0; // @[Mux.scala 19:72:@21629.4]
  assign _T_27694 = {conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,_T_27557}; // @[Mux.scala 19:72:@21644.4]
  assign _T_27696 = _T_2711 ? _T_27694 : 16'h0; // @[Mux.scala 19:72:@21645.4]
  assign _T_27711 = {conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,_T_27574}; // @[Mux.scala 19:72:@21660.4]
  assign _T_27713 = _T_2712 ? _T_27711 : 16'h0; // @[Mux.scala 19:72:@21661.4]
  assign _T_27714 = _T_27458 | _T_27475; // @[Mux.scala 19:72:@21662.4]
  assign _T_27715 = _T_27714 | _T_27492; // @[Mux.scala 19:72:@21663.4]
  assign _T_27716 = _T_27715 | _T_27509; // @[Mux.scala 19:72:@21664.4]
  assign _T_27717 = _T_27716 | _T_27526; // @[Mux.scala 19:72:@21665.4]
  assign _T_27718 = _T_27717 | _T_27543; // @[Mux.scala 19:72:@21666.4]
  assign _T_27719 = _T_27718 | _T_27560; // @[Mux.scala 19:72:@21667.4]
  assign _T_27720 = _T_27719 | _T_27577; // @[Mux.scala 19:72:@21668.4]
  assign _T_27721 = _T_27720 | _T_27594; // @[Mux.scala 19:72:@21669.4]
  assign _T_27722 = _T_27721 | _T_27611; // @[Mux.scala 19:72:@21670.4]
  assign _T_27723 = _T_27722 | _T_27628; // @[Mux.scala 19:72:@21671.4]
  assign _T_27724 = _T_27723 | _T_27645; // @[Mux.scala 19:72:@21672.4]
  assign _T_27725 = _T_27724 | _T_27662; // @[Mux.scala 19:72:@21673.4]
  assign _T_27726 = _T_27725 | _T_27679; // @[Mux.scala 19:72:@21674.4]
  assign _T_27727 = _T_27726 | _T_27696; // @[Mux.scala 19:72:@21675.4]
  assign _T_27728 = _T_27727 | _T_27713; // @[Mux.scala 19:72:@21676.4]
  assign _T_28306 = {conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0}; // @[Mux.scala 19:72:@22026.4]
  assign _T_28313 = {conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8}; // @[Mux.scala 19:72:@22033.4]
  assign _T_28314 = {conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,_T_28306}; // @[Mux.scala 19:72:@22034.4]
  assign _T_28316 = _T_2697 ? _T_28314 : 16'h0; // @[Mux.scala 19:72:@22035.4]
  assign _T_28323 = {conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1}; // @[Mux.scala 19:72:@22042.4]
  assign _T_28330 = {conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9}; // @[Mux.scala 19:72:@22049.4]
  assign _T_28331 = {conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,_T_28323}; // @[Mux.scala 19:72:@22050.4]
  assign _T_28333 = _T_2698 ? _T_28331 : 16'h0; // @[Mux.scala 19:72:@22051.4]
  assign _T_28340 = {conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2}; // @[Mux.scala 19:72:@22058.4]
  assign _T_28347 = {conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10}; // @[Mux.scala 19:72:@22065.4]
  assign _T_28348 = {conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,_T_28340}; // @[Mux.scala 19:72:@22066.4]
  assign _T_28350 = _T_2699 ? _T_28348 : 16'h0; // @[Mux.scala 19:72:@22067.4]
  assign _T_28357 = {conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3}; // @[Mux.scala 19:72:@22074.4]
  assign _T_28364 = {conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11}; // @[Mux.scala 19:72:@22081.4]
  assign _T_28365 = {conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,_T_28357}; // @[Mux.scala 19:72:@22082.4]
  assign _T_28367 = _T_2700 ? _T_28365 : 16'h0; // @[Mux.scala 19:72:@22083.4]
  assign _T_28374 = {conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4}; // @[Mux.scala 19:72:@22090.4]
  assign _T_28381 = {conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12}; // @[Mux.scala 19:72:@22097.4]
  assign _T_28382 = {conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,_T_28374}; // @[Mux.scala 19:72:@22098.4]
  assign _T_28384 = _T_2701 ? _T_28382 : 16'h0; // @[Mux.scala 19:72:@22099.4]
  assign _T_28391 = {conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5}; // @[Mux.scala 19:72:@22106.4]
  assign _T_28398 = {conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13}; // @[Mux.scala 19:72:@22113.4]
  assign _T_28399 = {conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,_T_28391}; // @[Mux.scala 19:72:@22114.4]
  assign _T_28401 = _T_2702 ? _T_28399 : 16'h0; // @[Mux.scala 19:72:@22115.4]
  assign _T_28408 = {conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6}; // @[Mux.scala 19:72:@22122.4]
  assign _T_28415 = {conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14}; // @[Mux.scala 19:72:@22129.4]
  assign _T_28416 = {conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,_T_28408}; // @[Mux.scala 19:72:@22130.4]
  assign _T_28418 = _T_2703 ? _T_28416 : 16'h0; // @[Mux.scala 19:72:@22131.4]
  assign _T_28425 = {conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7}; // @[Mux.scala 19:72:@22138.4]
  assign _T_28432 = {conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15}; // @[Mux.scala 19:72:@22145.4]
  assign _T_28433 = {conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,_T_28425}; // @[Mux.scala 19:72:@22146.4]
  assign _T_28435 = _T_2704 ? _T_28433 : 16'h0; // @[Mux.scala 19:72:@22147.4]
  assign _T_28450 = {conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,_T_28313}; // @[Mux.scala 19:72:@22162.4]
  assign _T_28452 = _T_2705 ? _T_28450 : 16'h0; // @[Mux.scala 19:72:@22163.4]
  assign _T_28467 = {conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,_T_28330}; // @[Mux.scala 19:72:@22178.4]
  assign _T_28469 = _T_2706 ? _T_28467 : 16'h0; // @[Mux.scala 19:72:@22179.4]
  assign _T_28484 = {conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,_T_28347}; // @[Mux.scala 19:72:@22194.4]
  assign _T_28486 = _T_2707 ? _T_28484 : 16'h0; // @[Mux.scala 19:72:@22195.4]
  assign _T_28501 = {conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,_T_28364}; // @[Mux.scala 19:72:@22210.4]
  assign _T_28503 = _T_2708 ? _T_28501 : 16'h0; // @[Mux.scala 19:72:@22211.4]
  assign _T_28518 = {conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,_T_28381}; // @[Mux.scala 19:72:@22226.4]
  assign _T_28520 = _T_2709 ? _T_28518 : 16'h0; // @[Mux.scala 19:72:@22227.4]
  assign _T_28535 = {conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,_T_28398}; // @[Mux.scala 19:72:@22242.4]
  assign _T_28537 = _T_2710 ? _T_28535 : 16'h0; // @[Mux.scala 19:72:@22243.4]
  assign _T_28552 = {conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,_T_28415}; // @[Mux.scala 19:72:@22258.4]
  assign _T_28554 = _T_2711 ? _T_28552 : 16'h0; // @[Mux.scala 19:72:@22259.4]
  assign _T_28569 = {conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,_T_28432}; // @[Mux.scala 19:72:@22274.4]
  assign _T_28571 = _T_2712 ? _T_28569 : 16'h0; // @[Mux.scala 19:72:@22275.4]
  assign _T_28572 = _T_28316 | _T_28333; // @[Mux.scala 19:72:@22276.4]
  assign _T_28573 = _T_28572 | _T_28350; // @[Mux.scala 19:72:@22277.4]
  assign _T_28574 = _T_28573 | _T_28367; // @[Mux.scala 19:72:@22278.4]
  assign _T_28575 = _T_28574 | _T_28384; // @[Mux.scala 19:72:@22279.4]
  assign _T_28576 = _T_28575 | _T_28401; // @[Mux.scala 19:72:@22280.4]
  assign _T_28577 = _T_28576 | _T_28418; // @[Mux.scala 19:72:@22281.4]
  assign _T_28578 = _T_28577 | _T_28435; // @[Mux.scala 19:72:@22282.4]
  assign _T_28579 = _T_28578 | _T_28452; // @[Mux.scala 19:72:@22283.4]
  assign _T_28580 = _T_28579 | _T_28469; // @[Mux.scala 19:72:@22284.4]
  assign _T_28581 = _T_28580 | _T_28486; // @[Mux.scala 19:72:@22285.4]
  assign _T_28582 = _T_28581 | _T_28503; // @[Mux.scala 19:72:@22286.4]
  assign _T_28583 = _T_28582 | _T_28520; // @[Mux.scala 19:72:@22287.4]
  assign _T_28584 = _T_28583 | _T_28537; // @[Mux.scala 19:72:@22288.4]
  assign _T_28585 = _T_28584 | _T_28554; // @[Mux.scala 19:72:@22289.4]
  assign _T_28586 = _T_28585 | _T_28571; // @[Mux.scala 19:72:@22290.4]
  assign _T_29164 = {conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0}; // @[Mux.scala 19:72:@22640.4]
  assign _T_29171 = {conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8}; // @[Mux.scala 19:72:@22647.4]
  assign _T_29172 = {conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,_T_29164}; // @[Mux.scala 19:72:@22648.4]
  assign _T_29174 = _T_2697 ? _T_29172 : 16'h0; // @[Mux.scala 19:72:@22649.4]
  assign _T_29181 = {conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1}; // @[Mux.scala 19:72:@22656.4]
  assign _T_29188 = {conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9}; // @[Mux.scala 19:72:@22663.4]
  assign _T_29189 = {conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,_T_29181}; // @[Mux.scala 19:72:@22664.4]
  assign _T_29191 = _T_2698 ? _T_29189 : 16'h0; // @[Mux.scala 19:72:@22665.4]
  assign _T_29198 = {conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2}; // @[Mux.scala 19:72:@22672.4]
  assign _T_29205 = {conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10}; // @[Mux.scala 19:72:@22679.4]
  assign _T_29206 = {conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,_T_29198}; // @[Mux.scala 19:72:@22680.4]
  assign _T_29208 = _T_2699 ? _T_29206 : 16'h0; // @[Mux.scala 19:72:@22681.4]
  assign _T_29215 = {conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3}; // @[Mux.scala 19:72:@22688.4]
  assign _T_29222 = {conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11}; // @[Mux.scala 19:72:@22695.4]
  assign _T_29223 = {conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,_T_29215}; // @[Mux.scala 19:72:@22696.4]
  assign _T_29225 = _T_2700 ? _T_29223 : 16'h0; // @[Mux.scala 19:72:@22697.4]
  assign _T_29232 = {conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4}; // @[Mux.scala 19:72:@22704.4]
  assign _T_29239 = {conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12}; // @[Mux.scala 19:72:@22711.4]
  assign _T_29240 = {conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,_T_29232}; // @[Mux.scala 19:72:@22712.4]
  assign _T_29242 = _T_2701 ? _T_29240 : 16'h0; // @[Mux.scala 19:72:@22713.4]
  assign _T_29249 = {conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5}; // @[Mux.scala 19:72:@22720.4]
  assign _T_29256 = {conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13}; // @[Mux.scala 19:72:@22727.4]
  assign _T_29257 = {conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,_T_29249}; // @[Mux.scala 19:72:@22728.4]
  assign _T_29259 = _T_2702 ? _T_29257 : 16'h0; // @[Mux.scala 19:72:@22729.4]
  assign _T_29266 = {conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6}; // @[Mux.scala 19:72:@22736.4]
  assign _T_29273 = {conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14}; // @[Mux.scala 19:72:@22743.4]
  assign _T_29274 = {conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,_T_29266}; // @[Mux.scala 19:72:@22744.4]
  assign _T_29276 = _T_2703 ? _T_29274 : 16'h0; // @[Mux.scala 19:72:@22745.4]
  assign _T_29283 = {conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7}; // @[Mux.scala 19:72:@22752.4]
  assign _T_29290 = {conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15}; // @[Mux.scala 19:72:@22759.4]
  assign _T_29291 = {conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,_T_29283}; // @[Mux.scala 19:72:@22760.4]
  assign _T_29293 = _T_2704 ? _T_29291 : 16'h0; // @[Mux.scala 19:72:@22761.4]
  assign _T_29308 = {conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,_T_29171}; // @[Mux.scala 19:72:@22776.4]
  assign _T_29310 = _T_2705 ? _T_29308 : 16'h0; // @[Mux.scala 19:72:@22777.4]
  assign _T_29325 = {conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,_T_29188}; // @[Mux.scala 19:72:@22792.4]
  assign _T_29327 = _T_2706 ? _T_29325 : 16'h0; // @[Mux.scala 19:72:@22793.4]
  assign _T_29342 = {conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,_T_29205}; // @[Mux.scala 19:72:@22808.4]
  assign _T_29344 = _T_2707 ? _T_29342 : 16'h0; // @[Mux.scala 19:72:@22809.4]
  assign _T_29359 = {conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,_T_29222}; // @[Mux.scala 19:72:@22824.4]
  assign _T_29361 = _T_2708 ? _T_29359 : 16'h0; // @[Mux.scala 19:72:@22825.4]
  assign _T_29376 = {conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,_T_29239}; // @[Mux.scala 19:72:@22840.4]
  assign _T_29378 = _T_2709 ? _T_29376 : 16'h0; // @[Mux.scala 19:72:@22841.4]
  assign _T_29393 = {conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,_T_29256}; // @[Mux.scala 19:72:@22856.4]
  assign _T_29395 = _T_2710 ? _T_29393 : 16'h0; // @[Mux.scala 19:72:@22857.4]
  assign _T_29410 = {conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,_T_29273}; // @[Mux.scala 19:72:@22872.4]
  assign _T_29412 = _T_2711 ? _T_29410 : 16'h0; // @[Mux.scala 19:72:@22873.4]
  assign _T_29427 = {conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,_T_29290}; // @[Mux.scala 19:72:@22888.4]
  assign _T_29429 = _T_2712 ? _T_29427 : 16'h0; // @[Mux.scala 19:72:@22889.4]
  assign _T_29430 = _T_29174 | _T_29191; // @[Mux.scala 19:72:@22890.4]
  assign _T_29431 = _T_29430 | _T_29208; // @[Mux.scala 19:72:@22891.4]
  assign _T_29432 = _T_29431 | _T_29225; // @[Mux.scala 19:72:@22892.4]
  assign _T_29433 = _T_29432 | _T_29242; // @[Mux.scala 19:72:@22893.4]
  assign _T_29434 = _T_29433 | _T_29259; // @[Mux.scala 19:72:@22894.4]
  assign _T_29435 = _T_29434 | _T_29276; // @[Mux.scala 19:72:@22895.4]
  assign _T_29436 = _T_29435 | _T_29293; // @[Mux.scala 19:72:@22896.4]
  assign _T_29437 = _T_29436 | _T_29310; // @[Mux.scala 19:72:@22897.4]
  assign _T_29438 = _T_29437 | _T_29327; // @[Mux.scala 19:72:@22898.4]
  assign _T_29439 = _T_29438 | _T_29344; // @[Mux.scala 19:72:@22899.4]
  assign _T_29440 = _T_29439 | _T_29361; // @[Mux.scala 19:72:@22900.4]
  assign _T_29441 = _T_29440 | _T_29378; // @[Mux.scala 19:72:@22901.4]
  assign _T_29442 = _T_29441 | _T_29395; // @[Mux.scala 19:72:@22902.4]
  assign _T_29443 = _T_29442 | _T_29412; // @[Mux.scala 19:72:@22903.4]
  assign _T_29444 = _T_29443 | _T_29429; // @[Mux.scala 19:72:@22904.4]
  assign _T_30022 = {conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0}; // @[Mux.scala 19:72:@23254.4]
  assign _T_30029 = {conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8}; // @[Mux.scala 19:72:@23261.4]
  assign _T_30030 = {conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,_T_30022}; // @[Mux.scala 19:72:@23262.4]
  assign _T_30032 = _T_2697 ? _T_30030 : 16'h0; // @[Mux.scala 19:72:@23263.4]
  assign _T_30039 = {conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1}; // @[Mux.scala 19:72:@23270.4]
  assign _T_30046 = {conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9}; // @[Mux.scala 19:72:@23277.4]
  assign _T_30047 = {conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,_T_30039}; // @[Mux.scala 19:72:@23278.4]
  assign _T_30049 = _T_2698 ? _T_30047 : 16'h0; // @[Mux.scala 19:72:@23279.4]
  assign _T_30056 = {conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2}; // @[Mux.scala 19:72:@23286.4]
  assign _T_30063 = {conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10}; // @[Mux.scala 19:72:@23293.4]
  assign _T_30064 = {conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,_T_30056}; // @[Mux.scala 19:72:@23294.4]
  assign _T_30066 = _T_2699 ? _T_30064 : 16'h0; // @[Mux.scala 19:72:@23295.4]
  assign _T_30073 = {conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3}; // @[Mux.scala 19:72:@23302.4]
  assign _T_30080 = {conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11}; // @[Mux.scala 19:72:@23309.4]
  assign _T_30081 = {conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,_T_30073}; // @[Mux.scala 19:72:@23310.4]
  assign _T_30083 = _T_2700 ? _T_30081 : 16'h0; // @[Mux.scala 19:72:@23311.4]
  assign _T_30090 = {conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4}; // @[Mux.scala 19:72:@23318.4]
  assign _T_30097 = {conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12}; // @[Mux.scala 19:72:@23325.4]
  assign _T_30098 = {conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,_T_30090}; // @[Mux.scala 19:72:@23326.4]
  assign _T_30100 = _T_2701 ? _T_30098 : 16'h0; // @[Mux.scala 19:72:@23327.4]
  assign _T_30107 = {conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5}; // @[Mux.scala 19:72:@23334.4]
  assign _T_30114 = {conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13}; // @[Mux.scala 19:72:@23341.4]
  assign _T_30115 = {conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,_T_30107}; // @[Mux.scala 19:72:@23342.4]
  assign _T_30117 = _T_2702 ? _T_30115 : 16'h0; // @[Mux.scala 19:72:@23343.4]
  assign _T_30124 = {conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6}; // @[Mux.scala 19:72:@23350.4]
  assign _T_30131 = {conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14}; // @[Mux.scala 19:72:@23357.4]
  assign _T_30132 = {conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,_T_30124}; // @[Mux.scala 19:72:@23358.4]
  assign _T_30134 = _T_2703 ? _T_30132 : 16'h0; // @[Mux.scala 19:72:@23359.4]
  assign _T_30141 = {conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7}; // @[Mux.scala 19:72:@23366.4]
  assign _T_30148 = {conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15}; // @[Mux.scala 19:72:@23373.4]
  assign _T_30149 = {conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,_T_30141}; // @[Mux.scala 19:72:@23374.4]
  assign _T_30151 = _T_2704 ? _T_30149 : 16'h0; // @[Mux.scala 19:72:@23375.4]
  assign _T_30166 = {conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,_T_30029}; // @[Mux.scala 19:72:@23390.4]
  assign _T_30168 = _T_2705 ? _T_30166 : 16'h0; // @[Mux.scala 19:72:@23391.4]
  assign _T_30183 = {conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,_T_30046}; // @[Mux.scala 19:72:@23406.4]
  assign _T_30185 = _T_2706 ? _T_30183 : 16'h0; // @[Mux.scala 19:72:@23407.4]
  assign _T_30200 = {conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,_T_30063}; // @[Mux.scala 19:72:@23422.4]
  assign _T_30202 = _T_2707 ? _T_30200 : 16'h0; // @[Mux.scala 19:72:@23423.4]
  assign _T_30217 = {conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,_T_30080}; // @[Mux.scala 19:72:@23438.4]
  assign _T_30219 = _T_2708 ? _T_30217 : 16'h0; // @[Mux.scala 19:72:@23439.4]
  assign _T_30234 = {conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,_T_30097}; // @[Mux.scala 19:72:@23454.4]
  assign _T_30236 = _T_2709 ? _T_30234 : 16'h0; // @[Mux.scala 19:72:@23455.4]
  assign _T_30251 = {conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,_T_30114}; // @[Mux.scala 19:72:@23470.4]
  assign _T_30253 = _T_2710 ? _T_30251 : 16'h0; // @[Mux.scala 19:72:@23471.4]
  assign _T_30268 = {conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,_T_30131}; // @[Mux.scala 19:72:@23486.4]
  assign _T_30270 = _T_2711 ? _T_30268 : 16'h0; // @[Mux.scala 19:72:@23487.4]
  assign _T_30285 = {conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,_T_30148}; // @[Mux.scala 19:72:@23502.4]
  assign _T_30287 = _T_2712 ? _T_30285 : 16'h0; // @[Mux.scala 19:72:@23503.4]
  assign _T_30288 = _T_30032 | _T_30049; // @[Mux.scala 19:72:@23504.4]
  assign _T_30289 = _T_30288 | _T_30066; // @[Mux.scala 19:72:@23505.4]
  assign _T_30290 = _T_30289 | _T_30083; // @[Mux.scala 19:72:@23506.4]
  assign _T_30291 = _T_30290 | _T_30100; // @[Mux.scala 19:72:@23507.4]
  assign _T_30292 = _T_30291 | _T_30117; // @[Mux.scala 19:72:@23508.4]
  assign _T_30293 = _T_30292 | _T_30134; // @[Mux.scala 19:72:@23509.4]
  assign _T_30294 = _T_30293 | _T_30151; // @[Mux.scala 19:72:@23510.4]
  assign _T_30295 = _T_30294 | _T_30168; // @[Mux.scala 19:72:@23511.4]
  assign _T_30296 = _T_30295 | _T_30185; // @[Mux.scala 19:72:@23512.4]
  assign _T_30297 = _T_30296 | _T_30202; // @[Mux.scala 19:72:@23513.4]
  assign _T_30298 = _T_30297 | _T_30219; // @[Mux.scala 19:72:@23514.4]
  assign _T_30299 = _T_30298 | _T_30236; // @[Mux.scala 19:72:@23515.4]
  assign _T_30300 = _T_30299 | _T_30253; // @[Mux.scala 19:72:@23516.4]
  assign _T_30301 = _T_30300 | _T_30270; // @[Mux.scala 19:72:@23517.4]
  assign _T_30302 = _T_30301 | _T_30287; // @[Mux.scala 19:72:@23518.4]
  assign _T_30880 = {conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0}; // @[Mux.scala 19:72:@23868.4]
  assign _T_30887 = {conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8}; // @[Mux.scala 19:72:@23875.4]
  assign _T_30888 = {conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,_T_30880}; // @[Mux.scala 19:72:@23876.4]
  assign _T_30890 = _T_2697 ? _T_30888 : 16'h0; // @[Mux.scala 19:72:@23877.4]
  assign _T_30897 = {conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1}; // @[Mux.scala 19:72:@23884.4]
  assign _T_30904 = {conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9}; // @[Mux.scala 19:72:@23891.4]
  assign _T_30905 = {conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,_T_30897}; // @[Mux.scala 19:72:@23892.4]
  assign _T_30907 = _T_2698 ? _T_30905 : 16'h0; // @[Mux.scala 19:72:@23893.4]
  assign _T_30914 = {conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2}; // @[Mux.scala 19:72:@23900.4]
  assign _T_30921 = {conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10}; // @[Mux.scala 19:72:@23907.4]
  assign _T_30922 = {conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,_T_30914}; // @[Mux.scala 19:72:@23908.4]
  assign _T_30924 = _T_2699 ? _T_30922 : 16'h0; // @[Mux.scala 19:72:@23909.4]
  assign _T_30931 = {conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3}; // @[Mux.scala 19:72:@23916.4]
  assign _T_30938 = {conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11}; // @[Mux.scala 19:72:@23923.4]
  assign _T_30939 = {conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,_T_30931}; // @[Mux.scala 19:72:@23924.4]
  assign _T_30941 = _T_2700 ? _T_30939 : 16'h0; // @[Mux.scala 19:72:@23925.4]
  assign _T_30948 = {conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4}; // @[Mux.scala 19:72:@23932.4]
  assign _T_30955 = {conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12}; // @[Mux.scala 19:72:@23939.4]
  assign _T_30956 = {conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,_T_30948}; // @[Mux.scala 19:72:@23940.4]
  assign _T_30958 = _T_2701 ? _T_30956 : 16'h0; // @[Mux.scala 19:72:@23941.4]
  assign _T_30965 = {conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5}; // @[Mux.scala 19:72:@23948.4]
  assign _T_30972 = {conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13}; // @[Mux.scala 19:72:@23955.4]
  assign _T_30973 = {conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,_T_30965}; // @[Mux.scala 19:72:@23956.4]
  assign _T_30975 = _T_2702 ? _T_30973 : 16'h0; // @[Mux.scala 19:72:@23957.4]
  assign _T_30982 = {conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6}; // @[Mux.scala 19:72:@23964.4]
  assign _T_30989 = {conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14}; // @[Mux.scala 19:72:@23971.4]
  assign _T_30990 = {conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,_T_30982}; // @[Mux.scala 19:72:@23972.4]
  assign _T_30992 = _T_2703 ? _T_30990 : 16'h0; // @[Mux.scala 19:72:@23973.4]
  assign _T_30999 = {conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7}; // @[Mux.scala 19:72:@23980.4]
  assign _T_31006 = {conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15}; // @[Mux.scala 19:72:@23987.4]
  assign _T_31007 = {conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,_T_30999}; // @[Mux.scala 19:72:@23988.4]
  assign _T_31009 = _T_2704 ? _T_31007 : 16'h0; // @[Mux.scala 19:72:@23989.4]
  assign _T_31024 = {conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,_T_30887}; // @[Mux.scala 19:72:@24004.4]
  assign _T_31026 = _T_2705 ? _T_31024 : 16'h0; // @[Mux.scala 19:72:@24005.4]
  assign _T_31041 = {conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,_T_30904}; // @[Mux.scala 19:72:@24020.4]
  assign _T_31043 = _T_2706 ? _T_31041 : 16'h0; // @[Mux.scala 19:72:@24021.4]
  assign _T_31058 = {conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,_T_30921}; // @[Mux.scala 19:72:@24036.4]
  assign _T_31060 = _T_2707 ? _T_31058 : 16'h0; // @[Mux.scala 19:72:@24037.4]
  assign _T_31075 = {conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,_T_30938}; // @[Mux.scala 19:72:@24052.4]
  assign _T_31077 = _T_2708 ? _T_31075 : 16'h0; // @[Mux.scala 19:72:@24053.4]
  assign _T_31092 = {conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,_T_30955}; // @[Mux.scala 19:72:@24068.4]
  assign _T_31094 = _T_2709 ? _T_31092 : 16'h0; // @[Mux.scala 19:72:@24069.4]
  assign _T_31109 = {conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,_T_30972}; // @[Mux.scala 19:72:@24084.4]
  assign _T_31111 = _T_2710 ? _T_31109 : 16'h0; // @[Mux.scala 19:72:@24085.4]
  assign _T_31126 = {conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,_T_30989}; // @[Mux.scala 19:72:@24100.4]
  assign _T_31128 = _T_2711 ? _T_31126 : 16'h0; // @[Mux.scala 19:72:@24101.4]
  assign _T_31143 = {conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,_T_31006}; // @[Mux.scala 19:72:@24116.4]
  assign _T_31145 = _T_2712 ? _T_31143 : 16'h0; // @[Mux.scala 19:72:@24117.4]
  assign _T_31146 = _T_30890 | _T_30907; // @[Mux.scala 19:72:@24118.4]
  assign _T_31147 = _T_31146 | _T_30924; // @[Mux.scala 19:72:@24119.4]
  assign _T_31148 = _T_31147 | _T_30941; // @[Mux.scala 19:72:@24120.4]
  assign _T_31149 = _T_31148 | _T_30958; // @[Mux.scala 19:72:@24121.4]
  assign _T_31150 = _T_31149 | _T_30975; // @[Mux.scala 19:72:@24122.4]
  assign _T_31151 = _T_31150 | _T_30992; // @[Mux.scala 19:72:@24123.4]
  assign _T_31152 = _T_31151 | _T_31009; // @[Mux.scala 19:72:@24124.4]
  assign _T_31153 = _T_31152 | _T_31026; // @[Mux.scala 19:72:@24125.4]
  assign _T_31154 = _T_31153 | _T_31043; // @[Mux.scala 19:72:@24126.4]
  assign _T_31155 = _T_31154 | _T_31060; // @[Mux.scala 19:72:@24127.4]
  assign _T_31156 = _T_31155 | _T_31077; // @[Mux.scala 19:72:@24128.4]
  assign _T_31157 = _T_31156 | _T_31094; // @[Mux.scala 19:72:@24129.4]
  assign _T_31158 = _T_31157 | _T_31111; // @[Mux.scala 19:72:@24130.4]
  assign _T_31159 = _T_31158 | _T_31128; // @[Mux.scala 19:72:@24131.4]
  assign _T_31160 = _T_31159 | _T_31145; // @[Mux.scala 19:72:@24132.4]
  assign _T_52334 = {storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0}; // @[Mux.scala 19:72:@24996.4]
  assign _T_52341 = {storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8}; // @[Mux.scala 19:72:@25003.4]
  assign _T_52342 = {storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,_T_52334}; // @[Mux.scala 19:72:@25004.4]
  assign _T_52344 = _T_2697 ? _T_52342 : 16'h0; // @[Mux.scala 19:72:@25005.4]
  assign _T_52351 = {storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1}; // @[Mux.scala 19:72:@25012.4]
  assign _T_52358 = {storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9}; // @[Mux.scala 19:72:@25019.4]
  assign _T_52359 = {storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,_T_52351}; // @[Mux.scala 19:72:@25020.4]
  assign _T_52361 = _T_2698 ? _T_52359 : 16'h0; // @[Mux.scala 19:72:@25021.4]
  assign _T_52368 = {storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2}; // @[Mux.scala 19:72:@25028.4]
  assign _T_52375 = {storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10}; // @[Mux.scala 19:72:@25035.4]
  assign _T_52376 = {storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,_T_52368}; // @[Mux.scala 19:72:@25036.4]
  assign _T_52378 = _T_2699 ? _T_52376 : 16'h0; // @[Mux.scala 19:72:@25037.4]
  assign _T_52385 = {storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3}; // @[Mux.scala 19:72:@25044.4]
  assign _T_52392 = {storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11}; // @[Mux.scala 19:72:@25051.4]
  assign _T_52393 = {storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,_T_52385}; // @[Mux.scala 19:72:@25052.4]
  assign _T_52395 = _T_2700 ? _T_52393 : 16'h0; // @[Mux.scala 19:72:@25053.4]
  assign _T_52402 = {storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4}; // @[Mux.scala 19:72:@25060.4]
  assign _T_52409 = {storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12}; // @[Mux.scala 19:72:@25067.4]
  assign _T_52410 = {storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,_T_52402}; // @[Mux.scala 19:72:@25068.4]
  assign _T_52412 = _T_2701 ? _T_52410 : 16'h0; // @[Mux.scala 19:72:@25069.4]
  assign _T_52419 = {storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5}; // @[Mux.scala 19:72:@25076.4]
  assign _T_52426 = {storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13}; // @[Mux.scala 19:72:@25083.4]
  assign _T_52427 = {storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,_T_52419}; // @[Mux.scala 19:72:@25084.4]
  assign _T_52429 = _T_2702 ? _T_52427 : 16'h0; // @[Mux.scala 19:72:@25085.4]
  assign _T_52436 = {storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6}; // @[Mux.scala 19:72:@25092.4]
  assign _T_52443 = {storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14}; // @[Mux.scala 19:72:@25099.4]
  assign _T_52444 = {storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,_T_52436}; // @[Mux.scala 19:72:@25100.4]
  assign _T_52446 = _T_2703 ? _T_52444 : 16'h0; // @[Mux.scala 19:72:@25101.4]
  assign _T_52453 = {storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7}; // @[Mux.scala 19:72:@25108.4]
  assign _T_52460 = {storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15}; // @[Mux.scala 19:72:@25115.4]
  assign _T_52461 = {storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,_T_52453}; // @[Mux.scala 19:72:@25116.4]
  assign _T_52463 = _T_2704 ? _T_52461 : 16'h0; // @[Mux.scala 19:72:@25117.4]
  assign _T_52478 = {storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,_T_52341}; // @[Mux.scala 19:72:@25132.4]
  assign _T_52480 = _T_2705 ? _T_52478 : 16'h0; // @[Mux.scala 19:72:@25133.4]
  assign _T_52495 = {storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,_T_52358}; // @[Mux.scala 19:72:@25148.4]
  assign _T_52497 = _T_2706 ? _T_52495 : 16'h0; // @[Mux.scala 19:72:@25149.4]
  assign _T_52512 = {storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,_T_52375}; // @[Mux.scala 19:72:@25164.4]
  assign _T_52514 = _T_2707 ? _T_52512 : 16'h0; // @[Mux.scala 19:72:@25165.4]
  assign _T_52529 = {storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,_T_52392}; // @[Mux.scala 19:72:@25180.4]
  assign _T_52531 = _T_2708 ? _T_52529 : 16'h0; // @[Mux.scala 19:72:@25181.4]
  assign _T_52546 = {storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,_T_52409}; // @[Mux.scala 19:72:@25196.4]
  assign _T_52548 = _T_2709 ? _T_52546 : 16'h0; // @[Mux.scala 19:72:@25197.4]
  assign _T_52563 = {storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,_T_52426}; // @[Mux.scala 19:72:@25212.4]
  assign _T_52565 = _T_2710 ? _T_52563 : 16'h0; // @[Mux.scala 19:72:@25213.4]
  assign _T_52580 = {storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,_T_52443}; // @[Mux.scala 19:72:@25228.4]
  assign _T_52582 = _T_2711 ? _T_52580 : 16'h0; // @[Mux.scala 19:72:@25229.4]
  assign _T_52597 = {storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,_T_52460}; // @[Mux.scala 19:72:@25244.4]
  assign _T_52599 = _T_2712 ? _T_52597 : 16'h0; // @[Mux.scala 19:72:@25245.4]
  assign _T_52600 = _T_52344 | _T_52361; // @[Mux.scala 19:72:@25246.4]
  assign _T_52601 = _T_52600 | _T_52378; // @[Mux.scala 19:72:@25247.4]
  assign _T_52602 = _T_52601 | _T_52395; // @[Mux.scala 19:72:@25248.4]
  assign _T_52603 = _T_52602 | _T_52412; // @[Mux.scala 19:72:@25249.4]
  assign _T_52604 = _T_52603 | _T_52429; // @[Mux.scala 19:72:@25250.4]
  assign _T_52605 = _T_52604 | _T_52446; // @[Mux.scala 19:72:@25251.4]
  assign _T_52606 = _T_52605 | _T_52463; // @[Mux.scala 19:72:@25252.4]
  assign _T_52607 = _T_52606 | _T_52480; // @[Mux.scala 19:72:@25253.4]
  assign _T_52608 = _T_52607 | _T_52497; // @[Mux.scala 19:72:@25254.4]
  assign _T_52609 = _T_52608 | _T_52514; // @[Mux.scala 19:72:@25255.4]
  assign _T_52610 = _T_52609 | _T_52531; // @[Mux.scala 19:72:@25256.4]
  assign _T_52611 = _T_52610 | _T_52548; // @[Mux.scala 19:72:@25257.4]
  assign _T_52612 = _T_52611 | _T_52565; // @[Mux.scala 19:72:@25258.4]
  assign _T_52613 = _T_52612 | _T_52582; // @[Mux.scala 19:72:@25259.4]
  assign _T_52614 = _T_52613 | _T_52599; // @[Mux.scala 19:72:@25260.4]
  assign _T_53192 = {storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0}; // @[Mux.scala 19:72:@25610.4]
  assign _T_53199 = {storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8}; // @[Mux.scala 19:72:@25617.4]
  assign _T_53200 = {storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,_T_53192}; // @[Mux.scala 19:72:@25618.4]
  assign _T_53202 = _T_2697 ? _T_53200 : 16'h0; // @[Mux.scala 19:72:@25619.4]
  assign _T_53209 = {storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1}; // @[Mux.scala 19:72:@25626.4]
  assign _T_53216 = {storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9}; // @[Mux.scala 19:72:@25633.4]
  assign _T_53217 = {storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,_T_53209}; // @[Mux.scala 19:72:@25634.4]
  assign _T_53219 = _T_2698 ? _T_53217 : 16'h0; // @[Mux.scala 19:72:@25635.4]
  assign _T_53226 = {storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2}; // @[Mux.scala 19:72:@25642.4]
  assign _T_53233 = {storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10}; // @[Mux.scala 19:72:@25649.4]
  assign _T_53234 = {storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,_T_53226}; // @[Mux.scala 19:72:@25650.4]
  assign _T_53236 = _T_2699 ? _T_53234 : 16'h0; // @[Mux.scala 19:72:@25651.4]
  assign _T_53243 = {storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3}; // @[Mux.scala 19:72:@25658.4]
  assign _T_53250 = {storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11}; // @[Mux.scala 19:72:@25665.4]
  assign _T_53251 = {storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,_T_53243}; // @[Mux.scala 19:72:@25666.4]
  assign _T_53253 = _T_2700 ? _T_53251 : 16'h0; // @[Mux.scala 19:72:@25667.4]
  assign _T_53260 = {storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4}; // @[Mux.scala 19:72:@25674.4]
  assign _T_53267 = {storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12}; // @[Mux.scala 19:72:@25681.4]
  assign _T_53268 = {storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,_T_53260}; // @[Mux.scala 19:72:@25682.4]
  assign _T_53270 = _T_2701 ? _T_53268 : 16'h0; // @[Mux.scala 19:72:@25683.4]
  assign _T_53277 = {storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5}; // @[Mux.scala 19:72:@25690.4]
  assign _T_53284 = {storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13}; // @[Mux.scala 19:72:@25697.4]
  assign _T_53285 = {storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,_T_53277}; // @[Mux.scala 19:72:@25698.4]
  assign _T_53287 = _T_2702 ? _T_53285 : 16'h0; // @[Mux.scala 19:72:@25699.4]
  assign _T_53294 = {storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6}; // @[Mux.scala 19:72:@25706.4]
  assign _T_53301 = {storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14}; // @[Mux.scala 19:72:@25713.4]
  assign _T_53302 = {storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,_T_53294}; // @[Mux.scala 19:72:@25714.4]
  assign _T_53304 = _T_2703 ? _T_53302 : 16'h0; // @[Mux.scala 19:72:@25715.4]
  assign _T_53311 = {storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7}; // @[Mux.scala 19:72:@25722.4]
  assign _T_53318 = {storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15}; // @[Mux.scala 19:72:@25729.4]
  assign _T_53319 = {storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,_T_53311}; // @[Mux.scala 19:72:@25730.4]
  assign _T_53321 = _T_2704 ? _T_53319 : 16'h0; // @[Mux.scala 19:72:@25731.4]
  assign _T_53336 = {storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,_T_53199}; // @[Mux.scala 19:72:@25746.4]
  assign _T_53338 = _T_2705 ? _T_53336 : 16'h0; // @[Mux.scala 19:72:@25747.4]
  assign _T_53353 = {storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,_T_53216}; // @[Mux.scala 19:72:@25762.4]
  assign _T_53355 = _T_2706 ? _T_53353 : 16'h0; // @[Mux.scala 19:72:@25763.4]
  assign _T_53370 = {storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,_T_53233}; // @[Mux.scala 19:72:@25778.4]
  assign _T_53372 = _T_2707 ? _T_53370 : 16'h0; // @[Mux.scala 19:72:@25779.4]
  assign _T_53387 = {storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,_T_53250}; // @[Mux.scala 19:72:@25794.4]
  assign _T_53389 = _T_2708 ? _T_53387 : 16'h0; // @[Mux.scala 19:72:@25795.4]
  assign _T_53404 = {storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,_T_53267}; // @[Mux.scala 19:72:@25810.4]
  assign _T_53406 = _T_2709 ? _T_53404 : 16'h0; // @[Mux.scala 19:72:@25811.4]
  assign _T_53421 = {storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,_T_53284}; // @[Mux.scala 19:72:@25826.4]
  assign _T_53423 = _T_2710 ? _T_53421 : 16'h0; // @[Mux.scala 19:72:@25827.4]
  assign _T_53438 = {storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,_T_53301}; // @[Mux.scala 19:72:@25842.4]
  assign _T_53440 = _T_2711 ? _T_53438 : 16'h0; // @[Mux.scala 19:72:@25843.4]
  assign _T_53455 = {storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,_T_53318}; // @[Mux.scala 19:72:@25858.4]
  assign _T_53457 = _T_2712 ? _T_53455 : 16'h0; // @[Mux.scala 19:72:@25859.4]
  assign _T_53458 = _T_53202 | _T_53219; // @[Mux.scala 19:72:@25860.4]
  assign _T_53459 = _T_53458 | _T_53236; // @[Mux.scala 19:72:@25861.4]
  assign _T_53460 = _T_53459 | _T_53253; // @[Mux.scala 19:72:@25862.4]
  assign _T_53461 = _T_53460 | _T_53270; // @[Mux.scala 19:72:@25863.4]
  assign _T_53462 = _T_53461 | _T_53287; // @[Mux.scala 19:72:@25864.4]
  assign _T_53463 = _T_53462 | _T_53304; // @[Mux.scala 19:72:@25865.4]
  assign _T_53464 = _T_53463 | _T_53321; // @[Mux.scala 19:72:@25866.4]
  assign _T_53465 = _T_53464 | _T_53338; // @[Mux.scala 19:72:@25867.4]
  assign _T_53466 = _T_53465 | _T_53355; // @[Mux.scala 19:72:@25868.4]
  assign _T_53467 = _T_53466 | _T_53372; // @[Mux.scala 19:72:@25869.4]
  assign _T_53468 = _T_53467 | _T_53389; // @[Mux.scala 19:72:@25870.4]
  assign _T_53469 = _T_53468 | _T_53406; // @[Mux.scala 19:72:@25871.4]
  assign _T_53470 = _T_53469 | _T_53423; // @[Mux.scala 19:72:@25872.4]
  assign _T_53471 = _T_53470 | _T_53440; // @[Mux.scala 19:72:@25873.4]
  assign _T_53472 = _T_53471 | _T_53457; // @[Mux.scala 19:72:@25874.4]
  assign _T_54050 = {storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0}; // @[Mux.scala 19:72:@26224.4]
  assign _T_54057 = {storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8}; // @[Mux.scala 19:72:@26231.4]
  assign _T_54058 = {storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,_T_54050}; // @[Mux.scala 19:72:@26232.4]
  assign _T_54060 = _T_2697 ? _T_54058 : 16'h0; // @[Mux.scala 19:72:@26233.4]
  assign _T_54067 = {storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1}; // @[Mux.scala 19:72:@26240.4]
  assign _T_54074 = {storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9}; // @[Mux.scala 19:72:@26247.4]
  assign _T_54075 = {storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,_T_54067}; // @[Mux.scala 19:72:@26248.4]
  assign _T_54077 = _T_2698 ? _T_54075 : 16'h0; // @[Mux.scala 19:72:@26249.4]
  assign _T_54084 = {storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2}; // @[Mux.scala 19:72:@26256.4]
  assign _T_54091 = {storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10}; // @[Mux.scala 19:72:@26263.4]
  assign _T_54092 = {storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,_T_54084}; // @[Mux.scala 19:72:@26264.4]
  assign _T_54094 = _T_2699 ? _T_54092 : 16'h0; // @[Mux.scala 19:72:@26265.4]
  assign _T_54101 = {storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3}; // @[Mux.scala 19:72:@26272.4]
  assign _T_54108 = {storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11}; // @[Mux.scala 19:72:@26279.4]
  assign _T_54109 = {storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,_T_54101}; // @[Mux.scala 19:72:@26280.4]
  assign _T_54111 = _T_2700 ? _T_54109 : 16'h0; // @[Mux.scala 19:72:@26281.4]
  assign _T_54118 = {storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4}; // @[Mux.scala 19:72:@26288.4]
  assign _T_54125 = {storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12}; // @[Mux.scala 19:72:@26295.4]
  assign _T_54126 = {storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,_T_54118}; // @[Mux.scala 19:72:@26296.4]
  assign _T_54128 = _T_2701 ? _T_54126 : 16'h0; // @[Mux.scala 19:72:@26297.4]
  assign _T_54135 = {storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5}; // @[Mux.scala 19:72:@26304.4]
  assign _T_54142 = {storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13}; // @[Mux.scala 19:72:@26311.4]
  assign _T_54143 = {storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,_T_54135}; // @[Mux.scala 19:72:@26312.4]
  assign _T_54145 = _T_2702 ? _T_54143 : 16'h0; // @[Mux.scala 19:72:@26313.4]
  assign _T_54152 = {storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6}; // @[Mux.scala 19:72:@26320.4]
  assign _T_54159 = {storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14}; // @[Mux.scala 19:72:@26327.4]
  assign _T_54160 = {storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,_T_54152}; // @[Mux.scala 19:72:@26328.4]
  assign _T_54162 = _T_2703 ? _T_54160 : 16'h0; // @[Mux.scala 19:72:@26329.4]
  assign _T_54169 = {storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7}; // @[Mux.scala 19:72:@26336.4]
  assign _T_54176 = {storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15}; // @[Mux.scala 19:72:@26343.4]
  assign _T_54177 = {storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,_T_54169}; // @[Mux.scala 19:72:@26344.4]
  assign _T_54179 = _T_2704 ? _T_54177 : 16'h0; // @[Mux.scala 19:72:@26345.4]
  assign _T_54194 = {storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,_T_54057}; // @[Mux.scala 19:72:@26360.4]
  assign _T_54196 = _T_2705 ? _T_54194 : 16'h0; // @[Mux.scala 19:72:@26361.4]
  assign _T_54211 = {storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,_T_54074}; // @[Mux.scala 19:72:@26376.4]
  assign _T_54213 = _T_2706 ? _T_54211 : 16'h0; // @[Mux.scala 19:72:@26377.4]
  assign _T_54228 = {storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,_T_54091}; // @[Mux.scala 19:72:@26392.4]
  assign _T_54230 = _T_2707 ? _T_54228 : 16'h0; // @[Mux.scala 19:72:@26393.4]
  assign _T_54245 = {storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,_T_54108}; // @[Mux.scala 19:72:@26408.4]
  assign _T_54247 = _T_2708 ? _T_54245 : 16'h0; // @[Mux.scala 19:72:@26409.4]
  assign _T_54262 = {storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,_T_54125}; // @[Mux.scala 19:72:@26424.4]
  assign _T_54264 = _T_2709 ? _T_54262 : 16'h0; // @[Mux.scala 19:72:@26425.4]
  assign _T_54279 = {storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,_T_54142}; // @[Mux.scala 19:72:@26440.4]
  assign _T_54281 = _T_2710 ? _T_54279 : 16'h0; // @[Mux.scala 19:72:@26441.4]
  assign _T_54296 = {storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,_T_54159}; // @[Mux.scala 19:72:@26456.4]
  assign _T_54298 = _T_2711 ? _T_54296 : 16'h0; // @[Mux.scala 19:72:@26457.4]
  assign _T_54313 = {storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,_T_54176}; // @[Mux.scala 19:72:@26472.4]
  assign _T_54315 = _T_2712 ? _T_54313 : 16'h0; // @[Mux.scala 19:72:@26473.4]
  assign _T_54316 = _T_54060 | _T_54077; // @[Mux.scala 19:72:@26474.4]
  assign _T_54317 = _T_54316 | _T_54094; // @[Mux.scala 19:72:@26475.4]
  assign _T_54318 = _T_54317 | _T_54111; // @[Mux.scala 19:72:@26476.4]
  assign _T_54319 = _T_54318 | _T_54128; // @[Mux.scala 19:72:@26477.4]
  assign _T_54320 = _T_54319 | _T_54145; // @[Mux.scala 19:72:@26478.4]
  assign _T_54321 = _T_54320 | _T_54162; // @[Mux.scala 19:72:@26479.4]
  assign _T_54322 = _T_54321 | _T_54179; // @[Mux.scala 19:72:@26480.4]
  assign _T_54323 = _T_54322 | _T_54196; // @[Mux.scala 19:72:@26481.4]
  assign _T_54324 = _T_54323 | _T_54213; // @[Mux.scala 19:72:@26482.4]
  assign _T_54325 = _T_54324 | _T_54230; // @[Mux.scala 19:72:@26483.4]
  assign _T_54326 = _T_54325 | _T_54247; // @[Mux.scala 19:72:@26484.4]
  assign _T_54327 = _T_54326 | _T_54264; // @[Mux.scala 19:72:@26485.4]
  assign _T_54328 = _T_54327 | _T_54281; // @[Mux.scala 19:72:@26486.4]
  assign _T_54329 = _T_54328 | _T_54298; // @[Mux.scala 19:72:@26487.4]
  assign _T_54330 = _T_54329 | _T_54315; // @[Mux.scala 19:72:@26488.4]
  assign _T_54908 = {storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0}; // @[Mux.scala 19:72:@26838.4]
  assign _T_54915 = {storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8}; // @[Mux.scala 19:72:@26845.4]
  assign _T_54916 = {storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,_T_54908}; // @[Mux.scala 19:72:@26846.4]
  assign _T_54918 = _T_2697 ? _T_54916 : 16'h0; // @[Mux.scala 19:72:@26847.4]
  assign _T_54925 = {storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1}; // @[Mux.scala 19:72:@26854.4]
  assign _T_54932 = {storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9}; // @[Mux.scala 19:72:@26861.4]
  assign _T_54933 = {storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,_T_54925}; // @[Mux.scala 19:72:@26862.4]
  assign _T_54935 = _T_2698 ? _T_54933 : 16'h0; // @[Mux.scala 19:72:@26863.4]
  assign _T_54942 = {storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2}; // @[Mux.scala 19:72:@26870.4]
  assign _T_54949 = {storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10}; // @[Mux.scala 19:72:@26877.4]
  assign _T_54950 = {storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,_T_54942}; // @[Mux.scala 19:72:@26878.4]
  assign _T_54952 = _T_2699 ? _T_54950 : 16'h0; // @[Mux.scala 19:72:@26879.4]
  assign _T_54959 = {storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3}; // @[Mux.scala 19:72:@26886.4]
  assign _T_54966 = {storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11}; // @[Mux.scala 19:72:@26893.4]
  assign _T_54967 = {storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,_T_54959}; // @[Mux.scala 19:72:@26894.4]
  assign _T_54969 = _T_2700 ? _T_54967 : 16'h0; // @[Mux.scala 19:72:@26895.4]
  assign _T_54976 = {storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4}; // @[Mux.scala 19:72:@26902.4]
  assign _T_54983 = {storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12}; // @[Mux.scala 19:72:@26909.4]
  assign _T_54984 = {storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,_T_54976}; // @[Mux.scala 19:72:@26910.4]
  assign _T_54986 = _T_2701 ? _T_54984 : 16'h0; // @[Mux.scala 19:72:@26911.4]
  assign _T_54993 = {storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5}; // @[Mux.scala 19:72:@26918.4]
  assign _T_55000 = {storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13}; // @[Mux.scala 19:72:@26925.4]
  assign _T_55001 = {storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,_T_54993}; // @[Mux.scala 19:72:@26926.4]
  assign _T_55003 = _T_2702 ? _T_55001 : 16'h0; // @[Mux.scala 19:72:@26927.4]
  assign _T_55010 = {storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6}; // @[Mux.scala 19:72:@26934.4]
  assign _T_55017 = {storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14}; // @[Mux.scala 19:72:@26941.4]
  assign _T_55018 = {storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,_T_55010}; // @[Mux.scala 19:72:@26942.4]
  assign _T_55020 = _T_2703 ? _T_55018 : 16'h0; // @[Mux.scala 19:72:@26943.4]
  assign _T_55027 = {storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7}; // @[Mux.scala 19:72:@26950.4]
  assign _T_55034 = {storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15}; // @[Mux.scala 19:72:@26957.4]
  assign _T_55035 = {storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,_T_55027}; // @[Mux.scala 19:72:@26958.4]
  assign _T_55037 = _T_2704 ? _T_55035 : 16'h0; // @[Mux.scala 19:72:@26959.4]
  assign _T_55052 = {storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,_T_54915}; // @[Mux.scala 19:72:@26974.4]
  assign _T_55054 = _T_2705 ? _T_55052 : 16'h0; // @[Mux.scala 19:72:@26975.4]
  assign _T_55069 = {storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,_T_54932}; // @[Mux.scala 19:72:@26990.4]
  assign _T_55071 = _T_2706 ? _T_55069 : 16'h0; // @[Mux.scala 19:72:@26991.4]
  assign _T_55086 = {storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,_T_54949}; // @[Mux.scala 19:72:@27006.4]
  assign _T_55088 = _T_2707 ? _T_55086 : 16'h0; // @[Mux.scala 19:72:@27007.4]
  assign _T_55103 = {storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,_T_54966}; // @[Mux.scala 19:72:@27022.4]
  assign _T_55105 = _T_2708 ? _T_55103 : 16'h0; // @[Mux.scala 19:72:@27023.4]
  assign _T_55120 = {storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,_T_54983}; // @[Mux.scala 19:72:@27038.4]
  assign _T_55122 = _T_2709 ? _T_55120 : 16'h0; // @[Mux.scala 19:72:@27039.4]
  assign _T_55137 = {storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,_T_55000}; // @[Mux.scala 19:72:@27054.4]
  assign _T_55139 = _T_2710 ? _T_55137 : 16'h0; // @[Mux.scala 19:72:@27055.4]
  assign _T_55154 = {storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,_T_55017}; // @[Mux.scala 19:72:@27070.4]
  assign _T_55156 = _T_2711 ? _T_55154 : 16'h0; // @[Mux.scala 19:72:@27071.4]
  assign _T_55171 = {storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,_T_55034}; // @[Mux.scala 19:72:@27086.4]
  assign _T_55173 = _T_2712 ? _T_55171 : 16'h0; // @[Mux.scala 19:72:@27087.4]
  assign _T_55174 = _T_54918 | _T_54935; // @[Mux.scala 19:72:@27088.4]
  assign _T_55175 = _T_55174 | _T_54952; // @[Mux.scala 19:72:@27089.4]
  assign _T_55176 = _T_55175 | _T_54969; // @[Mux.scala 19:72:@27090.4]
  assign _T_55177 = _T_55176 | _T_54986; // @[Mux.scala 19:72:@27091.4]
  assign _T_55178 = _T_55177 | _T_55003; // @[Mux.scala 19:72:@27092.4]
  assign _T_55179 = _T_55178 | _T_55020; // @[Mux.scala 19:72:@27093.4]
  assign _T_55180 = _T_55179 | _T_55037; // @[Mux.scala 19:72:@27094.4]
  assign _T_55181 = _T_55180 | _T_55054; // @[Mux.scala 19:72:@27095.4]
  assign _T_55182 = _T_55181 | _T_55071; // @[Mux.scala 19:72:@27096.4]
  assign _T_55183 = _T_55182 | _T_55088; // @[Mux.scala 19:72:@27097.4]
  assign _T_55184 = _T_55183 | _T_55105; // @[Mux.scala 19:72:@27098.4]
  assign _T_55185 = _T_55184 | _T_55122; // @[Mux.scala 19:72:@27099.4]
  assign _T_55186 = _T_55185 | _T_55139; // @[Mux.scala 19:72:@27100.4]
  assign _T_55187 = _T_55186 | _T_55156; // @[Mux.scala 19:72:@27101.4]
  assign _T_55188 = _T_55187 | _T_55173; // @[Mux.scala 19:72:@27102.4]
  assign _T_55766 = {storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0}; // @[Mux.scala 19:72:@27452.4]
  assign _T_55773 = {storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8}; // @[Mux.scala 19:72:@27459.4]
  assign _T_55774 = {storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,_T_55766}; // @[Mux.scala 19:72:@27460.4]
  assign _T_55776 = _T_2697 ? _T_55774 : 16'h0; // @[Mux.scala 19:72:@27461.4]
  assign _T_55783 = {storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1}; // @[Mux.scala 19:72:@27468.4]
  assign _T_55790 = {storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9}; // @[Mux.scala 19:72:@27475.4]
  assign _T_55791 = {storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,_T_55783}; // @[Mux.scala 19:72:@27476.4]
  assign _T_55793 = _T_2698 ? _T_55791 : 16'h0; // @[Mux.scala 19:72:@27477.4]
  assign _T_55800 = {storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2}; // @[Mux.scala 19:72:@27484.4]
  assign _T_55807 = {storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10}; // @[Mux.scala 19:72:@27491.4]
  assign _T_55808 = {storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,_T_55800}; // @[Mux.scala 19:72:@27492.4]
  assign _T_55810 = _T_2699 ? _T_55808 : 16'h0; // @[Mux.scala 19:72:@27493.4]
  assign _T_55817 = {storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3}; // @[Mux.scala 19:72:@27500.4]
  assign _T_55824 = {storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11}; // @[Mux.scala 19:72:@27507.4]
  assign _T_55825 = {storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,_T_55817}; // @[Mux.scala 19:72:@27508.4]
  assign _T_55827 = _T_2700 ? _T_55825 : 16'h0; // @[Mux.scala 19:72:@27509.4]
  assign _T_55834 = {storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4}; // @[Mux.scala 19:72:@27516.4]
  assign _T_55841 = {storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12}; // @[Mux.scala 19:72:@27523.4]
  assign _T_55842 = {storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,_T_55834}; // @[Mux.scala 19:72:@27524.4]
  assign _T_55844 = _T_2701 ? _T_55842 : 16'h0; // @[Mux.scala 19:72:@27525.4]
  assign _T_55851 = {storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5}; // @[Mux.scala 19:72:@27532.4]
  assign _T_55858 = {storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13}; // @[Mux.scala 19:72:@27539.4]
  assign _T_55859 = {storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,_T_55851}; // @[Mux.scala 19:72:@27540.4]
  assign _T_55861 = _T_2702 ? _T_55859 : 16'h0; // @[Mux.scala 19:72:@27541.4]
  assign _T_55868 = {storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6}; // @[Mux.scala 19:72:@27548.4]
  assign _T_55875 = {storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14}; // @[Mux.scala 19:72:@27555.4]
  assign _T_55876 = {storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,_T_55868}; // @[Mux.scala 19:72:@27556.4]
  assign _T_55878 = _T_2703 ? _T_55876 : 16'h0; // @[Mux.scala 19:72:@27557.4]
  assign _T_55885 = {storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7}; // @[Mux.scala 19:72:@27564.4]
  assign _T_55892 = {storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15}; // @[Mux.scala 19:72:@27571.4]
  assign _T_55893 = {storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,_T_55885}; // @[Mux.scala 19:72:@27572.4]
  assign _T_55895 = _T_2704 ? _T_55893 : 16'h0; // @[Mux.scala 19:72:@27573.4]
  assign _T_55910 = {storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,_T_55773}; // @[Mux.scala 19:72:@27588.4]
  assign _T_55912 = _T_2705 ? _T_55910 : 16'h0; // @[Mux.scala 19:72:@27589.4]
  assign _T_55927 = {storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,_T_55790}; // @[Mux.scala 19:72:@27604.4]
  assign _T_55929 = _T_2706 ? _T_55927 : 16'h0; // @[Mux.scala 19:72:@27605.4]
  assign _T_55944 = {storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,_T_55807}; // @[Mux.scala 19:72:@27620.4]
  assign _T_55946 = _T_2707 ? _T_55944 : 16'h0; // @[Mux.scala 19:72:@27621.4]
  assign _T_55961 = {storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,_T_55824}; // @[Mux.scala 19:72:@27636.4]
  assign _T_55963 = _T_2708 ? _T_55961 : 16'h0; // @[Mux.scala 19:72:@27637.4]
  assign _T_55978 = {storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,_T_55841}; // @[Mux.scala 19:72:@27652.4]
  assign _T_55980 = _T_2709 ? _T_55978 : 16'h0; // @[Mux.scala 19:72:@27653.4]
  assign _T_55995 = {storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,_T_55858}; // @[Mux.scala 19:72:@27668.4]
  assign _T_55997 = _T_2710 ? _T_55995 : 16'h0; // @[Mux.scala 19:72:@27669.4]
  assign _T_56012 = {storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,_T_55875}; // @[Mux.scala 19:72:@27684.4]
  assign _T_56014 = _T_2711 ? _T_56012 : 16'h0; // @[Mux.scala 19:72:@27685.4]
  assign _T_56029 = {storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,_T_55892}; // @[Mux.scala 19:72:@27700.4]
  assign _T_56031 = _T_2712 ? _T_56029 : 16'h0; // @[Mux.scala 19:72:@27701.4]
  assign _T_56032 = _T_55776 | _T_55793; // @[Mux.scala 19:72:@27702.4]
  assign _T_56033 = _T_56032 | _T_55810; // @[Mux.scala 19:72:@27703.4]
  assign _T_56034 = _T_56033 | _T_55827; // @[Mux.scala 19:72:@27704.4]
  assign _T_56035 = _T_56034 | _T_55844; // @[Mux.scala 19:72:@27705.4]
  assign _T_56036 = _T_56035 | _T_55861; // @[Mux.scala 19:72:@27706.4]
  assign _T_56037 = _T_56036 | _T_55878; // @[Mux.scala 19:72:@27707.4]
  assign _T_56038 = _T_56037 | _T_55895; // @[Mux.scala 19:72:@27708.4]
  assign _T_56039 = _T_56038 | _T_55912; // @[Mux.scala 19:72:@27709.4]
  assign _T_56040 = _T_56039 | _T_55929; // @[Mux.scala 19:72:@27710.4]
  assign _T_56041 = _T_56040 | _T_55946; // @[Mux.scala 19:72:@27711.4]
  assign _T_56042 = _T_56041 | _T_55963; // @[Mux.scala 19:72:@27712.4]
  assign _T_56043 = _T_56042 | _T_55980; // @[Mux.scala 19:72:@27713.4]
  assign _T_56044 = _T_56043 | _T_55997; // @[Mux.scala 19:72:@27714.4]
  assign _T_56045 = _T_56044 | _T_56014; // @[Mux.scala 19:72:@27715.4]
  assign _T_56046 = _T_56045 | _T_56031; // @[Mux.scala 19:72:@27716.4]
  assign _T_56624 = {storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0}; // @[Mux.scala 19:72:@28066.4]
  assign _T_56631 = {storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8}; // @[Mux.scala 19:72:@28073.4]
  assign _T_56632 = {storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,_T_56624}; // @[Mux.scala 19:72:@28074.4]
  assign _T_56634 = _T_2697 ? _T_56632 : 16'h0; // @[Mux.scala 19:72:@28075.4]
  assign _T_56641 = {storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1}; // @[Mux.scala 19:72:@28082.4]
  assign _T_56648 = {storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9}; // @[Mux.scala 19:72:@28089.4]
  assign _T_56649 = {storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,_T_56641}; // @[Mux.scala 19:72:@28090.4]
  assign _T_56651 = _T_2698 ? _T_56649 : 16'h0; // @[Mux.scala 19:72:@28091.4]
  assign _T_56658 = {storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2}; // @[Mux.scala 19:72:@28098.4]
  assign _T_56665 = {storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10}; // @[Mux.scala 19:72:@28105.4]
  assign _T_56666 = {storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,_T_56658}; // @[Mux.scala 19:72:@28106.4]
  assign _T_56668 = _T_2699 ? _T_56666 : 16'h0; // @[Mux.scala 19:72:@28107.4]
  assign _T_56675 = {storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3}; // @[Mux.scala 19:72:@28114.4]
  assign _T_56682 = {storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11}; // @[Mux.scala 19:72:@28121.4]
  assign _T_56683 = {storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,_T_56675}; // @[Mux.scala 19:72:@28122.4]
  assign _T_56685 = _T_2700 ? _T_56683 : 16'h0; // @[Mux.scala 19:72:@28123.4]
  assign _T_56692 = {storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4}; // @[Mux.scala 19:72:@28130.4]
  assign _T_56699 = {storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12}; // @[Mux.scala 19:72:@28137.4]
  assign _T_56700 = {storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,_T_56692}; // @[Mux.scala 19:72:@28138.4]
  assign _T_56702 = _T_2701 ? _T_56700 : 16'h0; // @[Mux.scala 19:72:@28139.4]
  assign _T_56709 = {storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5}; // @[Mux.scala 19:72:@28146.4]
  assign _T_56716 = {storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13}; // @[Mux.scala 19:72:@28153.4]
  assign _T_56717 = {storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,_T_56709}; // @[Mux.scala 19:72:@28154.4]
  assign _T_56719 = _T_2702 ? _T_56717 : 16'h0; // @[Mux.scala 19:72:@28155.4]
  assign _T_56726 = {storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6}; // @[Mux.scala 19:72:@28162.4]
  assign _T_56733 = {storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14}; // @[Mux.scala 19:72:@28169.4]
  assign _T_56734 = {storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,_T_56726}; // @[Mux.scala 19:72:@28170.4]
  assign _T_56736 = _T_2703 ? _T_56734 : 16'h0; // @[Mux.scala 19:72:@28171.4]
  assign _T_56743 = {storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7}; // @[Mux.scala 19:72:@28178.4]
  assign _T_56750 = {storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15}; // @[Mux.scala 19:72:@28185.4]
  assign _T_56751 = {storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,_T_56743}; // @[Mux.scala 19:72:@28186.4]
  assign _T_56753 = _T_2704 ? _T_56751 : 16'h0; // @[Mux.scala 19:72:@28187.4]
  assign _T_56768 = {storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,_T_56631}; // @[Mux.scala 19:72:@28202.4]
  assign _T_56770 = _T_2705 ? _T_56768 : 16'h0; // @[Mux.scala 19:72:@28203.4]
  assign _T_56785 = {storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,_T_56648}; // @[Mux.scala 19:72:@28218.4]
  assign _T_56787 = _T_2706 ? _T_56785 : 16'h0; // @[Mux.scala 19:72:@28219.4]
  assign _T_56802 = {storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,_T_56665}; // @[Mux.scala 19:72:@28234.4]
  assign _T_56804 = _T_2707 ? _T_56802 : 16'h0; // @[Mux.scala 19:72:@28235.4]
  assign _T_56819 = {storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,_T_56682}; // @[Mux.scala 19:72:@28250.4]
  assign _T_56821 = _T_2708 ? _T_56819 : 16'h0; // @[Mux.scala 19:72:@28251.4]
  assign _T_56836 = {storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,_T_56699}; // @[Mux.scala 19:72:@28266.4]
  assign _T_56838 = _T_2709 ? _T_56836 : 16'h0; // @[Mux.scala 19:72:@28267.4]
  assign _T_56853 = {storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,_T_56716}; // @[Mux.scala 19:72:@28282.4]
  assign _T_56855 = _T_2710 ? _T_56853 : 16'h0; // @[Mux.scala 19:72:@28283.4]
  assign _T_56870 = {storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,_T_56733}; // @[Mux.scala 19:72:@28298.4]
  assign _T_56872 = _T_2711 ? _T_56870 : 16'h0; // @[Mux.scala 19:72:@28299.4]
  assign _T_56887 = {storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,_T_56750}; // @[Mux.scala 19:72:@28314.4]
  assign _T_56889 = _T_2712 ? _T_56887 : 16'h0; // @[Mux.scala 19:72:@28315.4]
  assign _T_56890 = _T_56634 | _T_56651; // @[Mux.scala 19:72:@28316.4]
  assign _T_56891 = _T_56890 | _T_56668; // @[Mux.scala 19:72:@28317.4]
  assign _T_56892 = _T_56891 | _T_56685; // @[Mux.scala 19:72:@28318.4]
  assign _T_56893 = _T_56892 | _T_56702; // @[Mux.scala 19:72:@28319.4]
  assign _T_56894 = _T_56893 | _T_56719; // @[Mux.scala 19:72:@28320.4]
  assign _T_56895 = _T_56894 | _T_56736; // @[Mux.scala 19:72:@28321.4]
  assign _T_56896 = _T_56895 | _T_56753; // @[Mux.scala 19:72:@28322.4]
  assign _T_56897 = _T_56896 | _T_56770; // @[Mux.scala 19:72:@28323.4]
  assign _T_56898 = _T_56897 | _T_56787; // @[Mux.scala 19:72:@28324.4]
  assign _T_56899 = _T_56898 | _T_56804; // @[Mux.scala 19:72:@28325.4]
  assign _T_56900 = _T_56899 | _T_56821; // @[Mux.scala 19:72:@28326.4]
  assign _T_56901 = _T_56900 | _T_56838; // @[Mux.scala 19:72:@28327.4]
  assign _T_56902 = _T_56901 | _T_56855; // @[Mux.scala 19:72:@28328.4]
  assign _T_56903 = _T_56902 | _T_56872; // @[Mux.scala 19:72:@28329.4]
  assign _T_56904 = _T_56903 | _T_56889; // @[Mux.scala 19:72:@28330.4]
  assign _T_57482 = {storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0}; // @[Mux.scala 19:72:@28680.4]
  assign _T_57489 = {storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8}; // @[Mux.scala 19:72:@28687.4]
  assign _T_57490 = {storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,_T_57482}; // @[Mux.scala 19:72:@28688.4]
  assign _T_57492 = _T_2697 ? _T_57490 : 16'h0; // @[Mux.scala 19:72:@28689.4]
  assign _T_57499 = {storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1}; // @[Mux.scala 19:72:@28696.4]
  assign _T_57506 = {storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9}; // @[Mux.scala 19:72:@28703.4]
  assign _T_57507 = {storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,_T_57499}; // @[Mux.scala 19:72:@28704.4]
  assign _T_57509 = _T_2698 ? _T_57507 : 16'h0; // @[Mux.scala 19:72:@28705.4]
  assign _T_57516 = {storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2}; // @[Mux.scala 19:72:@28712.4]
  assign _T_57523 = {storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10}; // @[Mux.scala 19:72:@28719.4]
  assign _T_57524 = {storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,_T_57516}; // @[Mux.scala 19:72:@28720.4]
  assign _T_57526 = _T_2699 ? _T_57524 : 16'h0; // @[Mux.scala 19:72:@28721.4]
  assign _T_57533 = {storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3}; // @[Mux.scala 19:72:@28728.4]
  assign _T_57540 = {storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11}; // @[Mux.scala 19:72:@28735.4]
  assign _T_57541 = {storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,_T_57533}; // @[Mux.scala 19:72:@28736.4]
  assign _T_57543 = _T_2700 ? _T_57541 : 16'h0; // @[Mux.scala 19:72:@28737.4]
  assign _T_57550 = {storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4}; // @[Mux.scala 19:72:@28744.4]
  assign _T_57557 = {storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12}; // @[Mux.scala 19:72:@28751.4]
  assign _T_57558 = {storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,_T_57550}; // @[Mux.scala 19:72:@28752.4]
  assign _T_57560 = _T_2701 ? _T_57558 : 16'h0; // @[Mux.scala 19:72:@28753.4]
  assign _T_57567 = {storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5}; // @[Mux.scala 19:72:@28760.4]
  assign _T_57574 = {storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13}; // @[Mux.scala 19:72:@28767.4]
  assign _T_57575 = {storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,_T_57567}; // @[Mux.scala 19:72:@28768.4]
  assign _T_57577 = _T_2702 ? _T_57575 : 16'h0; // @[Mux.scala 19:72:@28769.4]
  assign _T_57584 = {storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6}; // @[Mux.scala 19:72:@28776.4]
  assign _T_57591 = {storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14}; // @[Mux.scala 19:72:@28783.4]
  assign _T_57592 = {storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,_T_57584}; // @[Mux.scala 19:72:@28784.4]
  assign _T_57594 = _T_2703 ? _T_57592 : 16'h0; // @[Mux.scala 19:72:@28785.4]
  assign _T_57601 = {storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7}; // @[Mux.scala 19:72:@28792.4]
  assign _T_57608 = {storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15}; // @[Mux.scala 19:72:@28799.4]
  assign _T_57609 = {storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,_T_57601}; // @[Mux.scala 19:72:@28800.4]
  assign _T_57611 = _T_2704 ? _T_57609 : 16'h0; // @[Mux.scala 19:72:@28801.4]
  assign _T_57626 = {storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,_T_57489}; // @[Mux.scala 19:72:@28816.4]
  assign _T_57628 = _T_2705 ? _T_57626 : 16'h0; // @[Mux.scala 19:72:@28817.4]
  assign _T_57643 = {storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,_T_57506}; // @[Mux.scala 19:72:@28832.4]
  assign _T_57645 = _T_2706 ? _T_57643 : 16'h0; // @[Mux.scala 19:72:@28833.4]
  assign _T_57660 = {storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,_T_57523}; // @[Mux.scala 19:72:@28848.4]
  assign _T_57662 = _T_2707 ? _T_57660 : 16'h0; // @[Mux.scala 19:72:@28849.4]
  assign _T_57677 = {storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,_T_57540}; // @[Mux.scala 19:72:@28864.4]
  assign _T_57679 = _T_2708 ? _T_57677 : 16'h0; // @[Mux.scala 19:72:@28865.4]
  assign _T_57694 = {storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,_T_57557}; // @[Mux.scala 19:72:@28880.4]
  assign _T_57696 = _T_2709 ? _T_57694 : 16'h0; // @[Mux.scala 19:72:@28881.4]
  assign _T_57711 = {storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,_T_57574}; // @[Mux.scala 19:72:@28896.4]
  assign _T_57713 = _T_2710 ? _T_57711 : 16'h0; // @[Mux.scala 19:72:@28897.4]
  assign _T_57728 = {storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,_T_57591}; // @[Mux.scala 19:72:@28912.4]
  assign _T_57730 = _T_2711 ? _T_57728 : 16'h0; // @[Mux.scala 19:72:@28913.4]
  assign _T_57745 = {storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,_T_57608}; // @[Mux.scala 19:72:@28928.4]
  assign _T_57747 = _T_2712 ? _T_57745 : 16'h0; // @[Mux.scala 19:72:@28929.4]
  assign _T_57748 = _T_57492 | _T_57509; // @[Mux.scala 19:72:@28930.4]
  assign _T_57749 = _T_57748 | _T_57526; // @[Mux.scala 19:72:@28931.4]
  assign _T_57750 = _T_57749 | _T_57543; // @[Mux.scala 19:72:@28932.4]
  assign _T_57751 = _T_57750 | _T_57560; // @[Mux.scala 19:72:@28933.4]
  assign _T_57752 = _T_57751 | _T_57577; // @[Mux.scala 19:72:@28934.4]
  assign _T_57753 = _T_57752 | _T_57594; // @[Mux.scala 19:72:@28935.4]
  assign _T_57754 = _T_57753 | _T_57611; // @[Mux.scala 19:72:@28936.4]
  assign _T_57755 = _T_57754 | _T_57628; // @[Mux.scala 19:72:@28937.4]
  assign _T_57756 = _T_57755 | _T_57645; // @[Mux.scala 19:72:@28938.4]
  assign _T_57757 = _T_57756 | _T_57662; // @[Mux.scala 19:72:@28939.4]
  assign _T_57758 = _T_57757 | _T_57679; // @[Mux.scala 19:72:@28940.4]
  assign _T_57759 = _T_57758 | _T_57696; // @[Mux.scala 19:72:@28941.4]
  assign _T_57760 = _T_57759 | _T_57713; // @[Mux.scala 19:72:@28942.4]
  assign _T_57761 = _T_57760 | _T_57730; // @[Mux.scala 19:72:@28943.4]
  assign _T_57762 = _T_57761 | _T_57747; // @[Mux.scala 19:72:@28944.4]
  assign _T_58340 = {storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0}; // @[Mux.scala 19:72:@29294.4]
  assign _T_58347 = {storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8}; // @[Mux.scala 19:72:@29301.4]
  assign _T_58348 = {storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,_T_58340}; // @[Mux.scala 19:72:@29302.4]
  assign _T_58350 = _T_2697 ? _T_58348 : 16'h0; // @[Mux.scala 19:72:@29303.4]
  assign _T_58357 = {storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1}; // @[Mux.scala 19:72:@29310.4]
  assign _T_58364 = {storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9}; // @[Mux.scala 19:72:@29317.4]
  assign _T_58365 = {storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,_T_58357}; // @[Mux.scala 19:72:@29318.4]
  assign _T_58367 = _T_2698 ? _T_58365 : 16'h0; // @[Mux.scala 19:72:@29319.4]
  assign _T_58374 = {storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2}; // @[Mux.scala 19:72:@29326.4]
  assign _T_58381 = {storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10}; // @[Mux.scala 19:72:@29333.4]
  assign _T_58382 = {storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,_T_58374}; // @[Mux.scala 19:72:@29334.4]
  assign _T_58384 = _T_2699 ? _T_58382 : 16'h0; // @[Mux.scala 19:72:@29335.4]
  assign _T_58391 = {storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3}; // @[Mux.scala 19:72:@29342.4]
  assign _T_58398 = {storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11}; // @[Mux.scala 19:72:@29349.4]
  assign _T_58399 = {storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,_T_58391}; // @[Mux.scala 19:72:@29350.4]
  assign _T_58401 = _T_2700 ? _T_58399 : 16'h0; // @[Mux.scala 19:72:@29351.4]
  assign _T_58408 = {storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4}; // @[Mux.scala 19:72:@29358.4]
  assign _T_58415 = {storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12}; // @[Mux.scala 19:72:@29365.4]
  assign _T_58416 = {storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,_T_58408}; // @[Mux.scala 19:72:@29366.4]
  assign _T_58418 = _T_2701 ? _T_58416 : 16'h0; // @[Mux.scala 19:72:@29367.4]
  assign _T_58425 = {storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5}; // @[Mux.scala 19:72:@29374.4]
  assign _T_58432 = {storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13}; // @[Mux.scala 19:72:@29381.4]
  assign _T_58433 = {storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,_T_58425}; // @[Mux.scala 19:72:@29382.4]
  assign _T_58435 = _T_2702 ? _T_58433 : 16'h0; // @[Mux.scala 19:72:@29383.4]
  assign _T_58442 = {storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6}; // @[Mux.scala 19:72:@29390.4]
  assign _T_58449 = {storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14}; // @[Mux.scala 19:72:@29397.4]
  assign _T_58450 = {storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,_T_58442}; // @[Mux.scala 19:72:@29398.4]
  assign _T_58452 = _T_2703 ? _T_58450 : 16'h0; // @[Mux.scala 19:72:@29399.4]
  assign _T_58459 = {storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7}; // @[Mux.scala 19:72:@29406.4]
  assign _T_58466 = {storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15}; // @[Mux.scala 19:72:@29413.4]
  assign _T_58467 = {storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,_T_58459}; // @[Mux.scala 19:72:@29414.4]
  assign _T_58469 = _T_2704 ? _T_58467 : 16'h0; // @[Mux.scala 19:72:@29415.4]
  assign _T_58484 = {storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,_T_58347}; // @[Mux.scala 19:72:@29430.4]
  assign _T_58486 = _T_2705 ? _T_58484 : 16'h0; // @[Mux.scala 19:72:@29431.4]
  assign _T_58501 = {storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,_T_58364}; // @[Mux.scala 19:72:@29446.4]
  assign _T_58503 = _T_2706 ? _T_58501 : 16'h0; // @[Mux.scala 19:72:@29447.4]
  assign _T_58518 = {storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,_T_58381}; // @[Mux.scala 19:72:@29462.4]
  assign _T_58520 = _T_2707 ? _T_58518 : 16'h0; // @[Mux.scala 19:72:@29463.4]
  assign _T_58535 = {storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,_T_58398}; // @[Mux.scala 19:72:@29478.4]
  assign _T_58537 = _T_2708 ? _T_58535 : 16'h0; // @[Mux.scala 19:72:@29479.4]
  assign _T_58552 = {storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,_T_58415}; // @[Mux.scala 19:72:@29494.4]
  assign _T_58554 = _T_2709 ? _T_58552 : 16'h0; // @[Mux.scala 19:72:@29495.4]
  assign _T_58569 = {storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,_T_58432}; // @[Mux.scala 19:72:@29510.4]
  assign _T_58571 = _T_2710 ? _T_58569 : 16'h0; // @[Mux.scala 19:72:@29511.4]
  assign _T_58586 = {storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,_T_58449}; // @[Mux.scala 19:72:@29526.4]
  assign _T_58588 = _T_2711 ? _T_58586 : 16'h0; // @[Mux.scala 19:72:@29527.4]
  assign _T_58603 = {storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,_T_58466}; // @[Mux.scala 19:72:@29542.4]
  assign _T_58605 = _T_2712 ? _T_58603 : 16'h0; // @[Mux.scala 19:72:@29543.4]
  assign _T_58606 = _T_58350 | _T_58367; // @[Mux.scala 19:72:@29544.4]
  assign _T_58607 = _T_58606 | _T_58384; // @[Mux.scala 19:72:@29545.4]
  assign _T_58608 = _T_58607 | _T_58401; // @[Mux.scala 19:72:@29546.4]
  assign _T_58609 = _T_58608 | _T_58418; // @[Mux.scala 19:72:@29547.4]
  assign _T_58610 = _T_58609 | _T_58435; // @[Mux.scala 19:72:@29548.4]
  assign _T_58611 = _T_58610 | _T_58452; // @[Mux.scala 19:72:@29549.4]
  assign _T_58612 = _T_58611 | _T_58469; // @[Mux.scala 19:72:@29550.4]
  assign _T_58613 = _T_58612 | _T_58486; // @[Mux.scala 19:72:@29551.4]
  assign _T_58614 = _T_58613 | _T_58503; // @[Mux.scala 19:72:@29552.4]
  assign _T_58615 = _T_58614 | _T_58520; // @[Mux.scala 19:72:@29553.4]
  assign _T_58616 = _T_58615 | _T_58537; // @[Mux.scala 19:72:@29554.4]
  assign _T_58617 = _T_58616 | _T_58554; // @[Mux.scala 19:72:@29555.4]
  assign _T_58618 = _T_58617 | _T_58571; // @[Mux.scala 19:72:@29556.4]
  assign _T_58619 = _T_58618 | _T_58588; // @[Mux.scala 19:72:@29557.4]
  assign _T_58620 = _T_58619 | _T_58605; // @[Mux.scala 19:72:@29558.4]
  assign _T_59198 = {storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0}; // @[Mux.scala 19:72:@29908.4]
  assign _T_59205 = {storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8}; // @[Mux.scala 19:72:@29915.4]
  assign _T_59206 = {storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,_T_59198}; // @[Mux.scala 19:72:@29916.4]
  assign _T_59208 = _T_2697 ? _T_59206 : 16'h0; // @[Mux.scala 19:72:@29917.4]
  assign _T_59215 = {storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1}; // @[Mux.scala 19:72:@29924.4]
  assign _T_59222 = {storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9}; // @[Mux.scala 19:72:@29931.4]
  assign _T_59223 = {storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,_T_59215}; // @[Mux.scala 19:72:@29932.4]
  assign _T_59225 = _T_2698 ? _T_59223 : 16'h0; // @[Mux.scala 19:72:@29933.4]
  assign _T_59232 = {storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2}; // @[Mux.scala 19:72:@29940.4]
  assign _T_59239 = {storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10}; // @[Mux.scala 19:72:@29947.4]
  assign _T_59240 = {storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,_T_59232}; // @[Mux.scala 19:72:@29948.4]
  assign _T_59242 = _T_2699 ? _T_59240 : 16'h0; // @[Mux.scala 19:72:@29949.4]
  assign _T_59249 = {storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3}; // @[Mux.scala 19:72:@29956.4]
  assign _T_59256 = {storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11}; // @[Mux.scala 19:72:@29963.4]
  assign _T_59257 = {storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,_T_59249}; // @[Mux.scala 19:72:@29964.4]
  assign _T_59259 = _T_2700 ? _T_59257 : 16'h0; // @[Mux.scala 19:72:@29965.4]
  assign _T_59266 = {storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4}; // @[Mux.scala 19:72:@29972.4]
  assign _T_59273 = {storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12}; // @[Mux.scala 19:72:@29979.4]
  assign _T_59274 = {storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,_T_59266}; // @[Mux.scala 19:72:@29980.4]
  assign _T_59276 = _T_2701 ? _T_59274 : 16'h0; // @[Mux.scala 19:72:@29981.4]
  assign _T_59283 = {storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5}; // @[Mux.scala 19:72:@29988.4]
  assign _T_59290 = {storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13}; // @[Mux.scala 19:72:@29995.4]
  assign _T_59291 = {storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,_T_59283}; // @[Mux.scala 19:72:@29996.4]
  assign _T_59293 = _T_2702 ? _T_59291 : 16'h0; // @[Mux.scala 19:72:@29997.4]
  assign _T_59300 = {storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6}; // @[Mux.scala 19:72:@30004.4]
  assign _T_59307 = {storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14}; // @[Mux.scala 19:72:@30011.4]
  assign _T_59308 = {storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,_T_59300}; // @[Mux.scala 19:72:@30012.4]
  assign _T_59310 = _T_2703 ? _T_59308 : 16'h0; // @[Mux.scala 19:72:@30013.4]
  assign _T_59317 = {storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7}; // @[Mux.scala 19:72:@30020.4]
  assign _T_59324 = {storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15}; // @[Mux.scala 19:72:@30027.4]
  assign _T_59325 = {storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,_T_59317}; // @[Mux.scala 19:72:@30028.4]
  assign _T_59327 = _T_2704 ? _T_59325 : 16'h0; // @[Mux.scala 19:72:@30029.4]
  assign _T_59342 = {storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,_T_59205}; // @[Mux.scala 19:72:@30044.4]
  assign _T_59344 = _T_2705 ? _T_59342 : 16'h0; // @[Mux.scala 19:72:@30045.4]
  assign _T_59359 = {storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,_T_59222}; // @[Mux.scala 19:72:@30060.4]
  assign _T_59361 = _T_2706 ? _T_59359 : 16'h0; // @[Mux.scala 19:72:@30061.4]
  assign _T_59376 = {storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,_T_59239}; // @[Mux.scala 19:72:@30076.4]
  assign _T_59378 = _T_2707 ? _T_59376 : 16'h0; // @[Mux.scala 19:72:@30077.4]
  assign _T_59393 = {storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,_T_59256}; // @[Mux.scala 19:72:@30092.4]
  assign _T_59395 = _T_2708 ? _T_59393 : 16'h0; // @[Mux.scala 19:72:@30093.4]
  assign _T_59410 = {storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,_T_59273}; // @[Mux.scala 19:72:@30108.4]
  assign _T_59412 = _T_2709 ? _T_59410 : 16'h0; // @[Mux.scala 19:72:@30109.4]
  assign _T_59427 = {storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,_T_59290}; // @[Mux.scala 19:72:@30124.4]
  assign _T_59429 = _T_2710 ? _T_59427 : 16'h0; // @[Mux.scala 19:72:@30125.4]
  assign _T_59444 = {storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,_T_59307}; // @[Mux.scala 19:72:@30140.4]
  assign _T_59446 = _T_2711 ? _T_59444 : 16'h0; // @[Mux.scala 19:72:@30141.4]
  assign _T_59461 = {storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,_T_59324}; // @[Mux.scala 19:72:@30156.4]
  assign _T_59463 = _T_2712 ? _T_59461 : 16'h0; // @[Mux.scala 19:72:@30157.4]
  assign _T_59464 = _T_59208 | _T_59225; // @[Mux.scala 19:72:@30158.4]
  assign _T_59465 = _T_59464 | _T_59242; // @[Mux.scala 19:72:@30159.4]
  assign _T_59466 = _T_59465 | _T_59259; // @[Mux.scala 19:72:@30160.4]
  assign _T_59467 = _T_59466 | _T_59276; // @[Mux.scala 19:72:@30161.4]
  assign _T_59468 = _T_59467 | _T_59293; // @[Mux.scala 19:72:@30162.4]
  assign _T_59469 = _T_59468 | _T_59310; // @[Mux.scala 19:72:@30163.4]
  assign _T_59470 = _T_59469 | _T_59327; // @[Mux.scala 19:72:@30164.4]
  assign _T_59471 = _T_59470 | _T_59344; // @[Mux.scala 19:72:@30165.4]
  assign _T_59472 = _T_59471 | _T_59361; // @[Mux.scala 19:72:@30166.4]
  assign _T_59473 = _T_59472 | _T_59378; // @[Mux.scala 19:72:@30167.4]
  assign _T_59474 = _T_59473 | _T_59395; // @[Mux.scala 19:72:@30168.4]
  assign _T_59475 = _T_59474 | _T_59412; // @[Mux.scala 19:72:@30169.4]
  assign _T_59476 = _T_59475 | _T_59429; // @[Mux.scala 19:72:@30170.4]
  assign _T_59477 = _T_59476 | _T_59446; // @[Mux.scala 19:72:@30171.4]
  assign _T_59478 = _T_59477 | _T_59463; // @[Mux.scala 19:72:@30172.4]
  assign _T_60056 = {storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0}; // @[Mux.scala 19:72:@30522.4]
  assign _T_60063 = {storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8}; // @[Mux.scala 19:72:@30529.4]
  assign _T_60064 = {storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,_T_60056}; // @[Mux.scala 19:72:@30530.4]
  assign _T_60066 = _T_2697 ? _T_60064 : 16'h0; // @[Mux.scala 19:72:@30531.4]
  assign _T_60073 = {storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1}; // @[Mux.scala 19:72:@30538.4]
  assign _T_60080 = {storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9}; // @[Mux.scala 19:72:@30545.4]
  assign _T_60081 = {storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,_T_60073}; // @[Mux.scala 19:72:@30546.4]
  assign _T_60083 = _T_2698 ? _T_60081 : 16'h0; // @[Mux.scala 19:72:@30547.4]
  assign _T_60090 = {storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2}; // @[Mux.scala 19:72:@30554.4]
  assign _T_60097 = {storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10}; // @[Mux.scala 19:72:@30561.4]
  assign _T_60098 = {storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,_T_60090}; // @[Mux.scala 19:72:@30562.4]
  assign _T_60100 = _T_2699 ? _T_60098 : 16'h0; // @[Mux.scala 19:72:@30563.4]
  assign _T_60107 = {storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3}; // @[Mux.scala 19:72:@30570.4]
  assign _T_60114 = {storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11}; // @[Mux.scala 19:72:@30577.4]
  assign _T_60115 = {storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,_T_60107}; // @[Mux.scala 19:72:@30578.4]
  assign _T_60117 = _T_2700 ? _T_60115 : 16'h0; // @[Mux.scala 19:72:@30579.4]
  assign _T_60124 = {storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4}; // @[Mux.scala 19:72:@30586.4]
  assign _T_60131 = {storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12}; // @[Mux.scala 19:72:@30593.4]
  assign _T_60132 = {storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,_T_60124}; // @[Mux.scala 19:72:@30594.4]
  assign _T_60134 = _T_2701 ? _T_60132 : 16'h0; // @[Mux.scala 19:72:@30595.4]
  assign _T_60141 = {storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5}; // @[Mux.scala 19:72:@30602.4]
  assign _T_60148 = {storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13}; // @[Mux.scala 19:72:@30609.4]
  assign _T_60149 = {storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,_T_60141}; // @[Mux.scala 19:72:@30610.4]
  assign _T_60151 = _T_2702 ? _T_60149 : 16'h0; // @[Mux.scala 19:72:@30611.4]
  assign _T_60158 = {storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6}; // @[Mux.scala 19:72:@30618.4]
  assign _T_60165 = {storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14}; // @[Mux.scala 19:72:@30625.4]
  assign _T_60166 = {storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,_T_60158}; // @[Mux.scala 19:72:@30626.4]
  assign _T_60168 = _T_2703 ? _T_60166 : 16'h0; // @[Mux.scala 19:72:@30627.4]
  assign _T_60175 = {storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7}; // @[Mux.scala 19:72:@30634.4]
  assign _T_60182 = {storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15}; // @[Mux.scala 19:72:@30641.4]
  assign _T_60183 = {storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,_T_60175}; // @[Mux.scala 19:72:@30642.4]
  assign _T_60185 = _T_2704 ? _T_60183 : 16'h0; // @[Mux.scala 19:72:@30643.4]
  assign _T_60200 = {storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,_T_60063}; // @[Mux.scala 19:72:@30658.4]
  assign _T_60202 = _T_2705 ? _T_60200 : 16'h0; // @[Mux.scala 19:72:@30659.4]
  assign _T_60217 = {storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,_T_60080}; // @[Mux.scala 19:72:@30674.4]
  assign _T_60219 = _T_2706 ? _T_60217 : 16'h0; // @[Mux.scala 19:72:@30675.4]
  assign _T_60234 = {storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,_T_60097}; // @[Mux.scala 19:72:@30690.4]
  assign _T_60236 = _T_2707 ? _T_60234 : 16'h0; // @[Mux.scala 19:72:@30691.4]
  assign _T_60251 = {storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,_T_60114}; // @[Mux.scala 19:72:@30706.4]
  assign _T_60253 = _T_2708 ? _T_60251 : 16'h0; // @[Mux.scala 19:72:@30707.4]
  assign _T_60268 = {storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,_T_60131}; // @[Mux.scala 19:72:@30722.4]
  assign _T_60270 = _T_2709 ? _T_60268 : 16'h0; // @[Mux.scala 19:72:@30723.4]
  assign _T_60285 = {storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,_T_60148}; // @[Mux.scala 19:72:@30738.4]
  assign _T_60287 = _T_2710 ? _T_60285 : 16'h0; // @[Mux.scala 19:72:@30739.4]
  assign _T_60302 = {storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,_T_60165}; // @[Mux.scala 19:72:@30754.4]
  assign _T_60304 = _T_2711 ? _T_60302 : 16'h0; // @[Mux.scala 19:72:@30755.4]
  assign _T_60319 = {storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,_T_60182}; // @[Mux.scala 19:72:@30770.4]
  assign _T_60321 = _T_2712 ? _T_60319 : 16'h0; // @[Mux.scala 19:72:@30771.4]
  assign _T_60322 = _T_60066 | _T_60083; // @[Mux.scala 19:72:@30772.4]
  assign _T_60323 = _T_60322 | _T_60100; // @[Mux.scala 19:72:@30773.4]
  assign _T_60324 = _T_60323 | _T_60117; // @[Mux.scala 19:72:@30774.4]
  assign _T_60325 = _T_60324 | _T_60134; // @[Mux.scala 19:72:@30775.4]
  assign _T_60326 = _T_60325 | _T_60151; // @[Mux.scala 19:72:@30776.4]
  assign _T_60327 = _T_60326 | _T_60168; // @[Mux.scala 19:72:@30777.4]
  assign _T_60328 = _T_60327 | _T_60185; // @[Mux.scala 19:72:@30778.4]
  assign _T_60329 = _T_60328 | _T_60202; // @[Mux.scala 19:72:@30779.4]
  assign _T_60330 = _T_60329 | _T_60219; // @[Mux.scala 19:72:@30780.4]
  assign _T_60331 = _T_60330 | _T_60236; // @[Mux.scala 19:72:@30781.4]
  assign _T_60332 = _T_60331 | _T_60253; // @[Mux.scala 19:72:@30782.4]
  assign _T_60333 = _T_60332 | _T_60270; // @[Mux.scala 19:72:@30783.4]
  assign _T_60334 = _T_60333 | _T_60287; // @[Mux.scala 19:72:@30784.4]
  assign _T_60335 = _T_60334 | _T_60304; // @[Mux.scala 19:72:@30785.4]
  assign _T_60336 = _T_60335 | _T_60321; // @[Mux.scala 19:72:@30786.4]
  assign _T_60914 = {storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0}; // @[Mux.scala 19:72:@31136.4]
  assign _T_60921 = {storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8}; // @[Mux.scala 19:72:@31143.4]
  assign _T_60922 = {storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,_T_60914}; // @[Mux.scala 19:72:@31144.4]
  assign _T_60924 = _T_2697 ? _T_60922 : 16'h0; // @[Mux.scala 19:72:@31145.4]
  assign _T_60931 = {storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1}; // @[Mux.scala 19:72:@31152.4]
  assign _T_60938 = {storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9}; // @[Mux.scala 19:72:@31159.4]
  assign _T_60939 = {storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,_T_60931}; // @[Mux.scala 19:72:@31160.4]
  assign _T_60941 = _T_2698 ? _T_60939 : 16'h0; // @[Mux.scala 19:72:@31161.4]
  assign _T_60948 = {storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2}; // @[Mux.scala 19:72:@31168.4]
  assign _T_60955 = {storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10}; // @[Mux.scala 19:72:@31175.4]
  assign _T_60956 = {storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,_T_60948}; // @[Mux.scala 19:72:@31176.4]
  assign _T_60958 = _T_2699 ? _T_60956 : 16'h0; // @[Mux.scala 19:72:@31177.4]
  assign _T_60965 = {storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3}; // @[Mux.scala 19:72:@31184.4]
  assign _T_60972 = {storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11}; // @[Mux.scala 19:72:@31191.4]
  assign _T_60973 = {storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,_T_60965}; // @[Mux.scala 19:72:@31192.4]
  assign _T_60975 = _T_2700 ? _T_60973 : 16'h0; // @[Mux.scala 19:72:@31193.4]
  assign _T_60982 = {storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4}; // @[Mux.scala 19:72:@31200.4]
  assign _T_60989 = {storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12}; // @[Mux.scala 19:72:@31207.4]
  assign _T_60990 = {storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,_T_60982}; // @[Mux.scala 19:72:@31208.4]
  assign _T_60992 = _T_2701 ? _T_60990 : 16'h0; // @[Mux.scala 19:72:@31209.4]
  assign _T_60999 = {storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5}; // @[Mux.scala 19:72:@31216.4]
  assign _T_61006 = {storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13}; // @[Mux.scala 19:72:@31223.4]
  assign _T_61007 = {storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,_T_60999}; // @[Mux.scala 19:72:@31224.4]
  assign _T_61009 = _T_2702 ? _T_61007 : 16'h0; // @[Mux.scala 19:72:@31225.4]
  assign _T_61016 = {storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6}; // @[Mux.scala 19:72:@31232.4]
  assign _T_61023 = {storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14}; // @[Mux.scala 19:72:@31239.4]
  assign _T_61024 = {storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,_T_61016}; // @[Mux.scala 19:72:@31240.4]
  assign _T_61026 = _T_2703 ? _T_61024 : 16'h0; // @[Mux.scala 19:72:@31241.4]
  assign _T_61033 = {storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7}; // @[Mux.scala 19:72:@31248.4]
  assign _T_61040 = {storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15}; // @[Mux.scala 19:72:@31255.4]
  assign _T_61041 = {storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,_T_61033}; // @[Mux.scala 19:72:@31256.4]
  assign _T_61043 = _T_2704 ? _T_61041 : 16'h0; // @[Mux.scala 19:72:@31257.4]
  assign _T_61058 = {storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,_T_60921}; // @[Mux.scala 19:72:@31272.4]
  assign _T_61060 = _T_2705 ? _T_61058 : 16'h0; // @[Mux.scala 19:72:@31273.4]
  assign _T_61075 = {storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,_T_60938}; // @[Mux.scala 19:72:@31288.4]
  assign _T_61077 = _T_2706 ? _T_61075 : 16'h0; // @[Mux.scala 19:72:@31289.4]
  assign _T_61092 = {storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,_T_60955}; // @[Mux.scala 19:72:@31304.4]
  assign _T_61094 = _T_2707 ? _T_61092 : 16'h0; // @[Mux.scala 19:72:@31305.4]
  assign _T_61109 = {storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,_T_60972}; // @[Mux.scala 19:72:@31320.4]
  assign _T_61111 = _T_2708 ? _T_61109 : 16'h0; // @[Mux.scala 19:72:@31321.4]
  assign _T_61126 = {storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,_T_60989}; // @[Mux.scala 19:72:@31336.4]
  assign _T_61128 = _T_2709 ? _T_61126 : 16'h0; // @[Mux.scala 19:72:@31337.4]
  assign _T_61143 = {storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,_T_61006}; // @[Mux.scala 19:72:@31352.4]
  assign _T_61145 = _T_2710 ? _T_61143 : 16'h0; // @[Mux.scala 19:72:@31353.4]
  assign _T_61160 = {storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,_T_61023}; // @[Mux.scala 19:72:@31368.4]
  assign _T_61162 = _T_2711 ? _T_61160 : 16'h0; // @[Mux.scala 19:72:@31369.4]
  assign _T_61177 = {storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,_T_61040}; // @[Mux.scala 19:72:@31384.4]
  assign _T_61179 = _T_2712 ? _T_61177 : 16'h0; // @[Mux.scala 19:72:@31385.4]
  assign _T_61180 = _T_60924 | _T_60941; // @[Mux.scala 19:72:@31386.4]
  assign _T_61181 = _T_61180 | _T_60958; // @[Mux.scala 19:72:@31387.4]
  assign _T_61182 = _T_61181 | _T_60975; // @[Mux.scala 19:72:@31388.4]
  assign _T_61183 = _T_61182 | _T_60992; // @[Mux.scala 19:72:@31389.4]
  assign _T_61184 = _T_61183 | _T_61009; // @[Mux.scala 19:72:@31390.4]
  assign _T_61185 = _T_61184 | _T_61026; // @[Mux.scala 19:72:@31391.4]
  assign _T_61186 = _T_61185 | _T_61043; // @[Mux.scala 19:72:@31392.4]
  assign _T_61187 = _T_61186 | _T_61060; // @[Mux.scala 19:72:@31393.4]
  assign _T_61188 = _T_61187 | _T_61077; // @[Mux.scala 19:72:@31394.4]
  assign _T_61189 = _T_61188 | _T_61094; // @[Mux.scala 19:72:@31395.4]
  assign _T_61190 = _T_61189 | _T_61111; // @[Mux.scala 19:72:@31396.4]
  assign _T_61191 = _T_61190 | _T_61128; // @[Mux.scala 19:72:@31397.4]
  assign _T_61192 = _T_61191 | _T_61145; // @[Mux.scala 19:72:@31398.4]
  assign _T_61193 = _T_61192 | _T_61162; // @[Mux.scala 19:72:@31399.4]
  assign _T_61194 = _T_61193 | _T_61179; // @[Mux.scala 19:72:@31400.4]
  assign _T_61772 = {storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0}; // @[Mux.scala 19:72:@31750.4]
  assign _T_61779 = {storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8}; // @[Mux.scala 19:72:@31757.4]
  assign _T_61780 = {storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,_T_61772}; // @[Mux.scala 19:72:@31758.4]
  assign _T_61782 = _T_2697 ? _T_61780 : 16'h0; // @[Mux.scala 19:72:@31759.4]
  assign _T_61789 = {storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1}; // @[Mux.scala 19:72:@31766.4]
  assign _T_61796 = {storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9}; // @[Mux.scala 19:72:@31773.4]
  assign _T_61797 = {storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,_T_61789}; // @[Mux.scala 19:72:@31774.4]
  assign _T_61799 = _T_2698 ? _T_61797 : 16'h0; // @[Mux.scala 19:72:@31775.4]
  assign _T_61806 = {storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2}; // @[Mux.scala 19:72:@31782.4]
  assign _T_61813 = {storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10}; // @[Mux.scala 19:72:@31789.4]
  assign _T_61814 = {storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,_T_61806}; // @[Mux.scala 19:72:@31790.4]
  assign _T_61816 = _T_2699 ? _T_61814 : 16'h0; // @[Mux.scala 19:72:@31791.4]
  assign _T_61823 = {storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3}; // @[Mux.scala 19:72:@31798.4]
  assign _T_61830 = {storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11}; // @[Mux.scala 19:72:@31805.4]
  assign _T_61831 = {storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,_T_61823}; // @[Mux.scala 19:72:@31806.4]
  assign _T_61833 = _T_2700 ? _T_61831 : 16'h0; // @[Mux.scala 19:72:@31807.4]
  assign _T_61840 = {storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4}; // @[Mux.scala 19:72:@31814.4]
  assign _T_61847 = {storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12}; // @[Mux.scala 19:72:@31821.4]
  assign _T_61848 = {storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,_T_61840}; // @[Mux.scala 19:72:@31822.4]
  assign _T_61850 = _T_2701 ? _T_61848 : 16'h0; // @[Mux.scala 19:72:@31823.4]
  assign _T_61857 = {storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5}; // @[Mux.scala 19:72:@31830.4]
  assign _T_61864 = {storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13}; // @[Mux.scala 19:72:@31837.4]
  assign _T_61865 = {storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,_T_61857}; // @[Mux.scala 19:72:@31838.4]
  assign _T_61867 = _T_2702 ? _T_61865 : 16'h0; // @[Mux.scala 19:72:@31839.4]
  assign _T_61874 = {storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6}; // @[Mux.scala 19:72:@31846.4]
  assign _T_61881 = {storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14}; // @[Mux.scala 19:72:@31853.4]
  assign _T_61882 = {storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,_T_61874}; // @[Mux.scala 19:72:@31854.4]
  assign _T_61884 = _T_2703 ? _T_61882 : 16'h0; // @[Mux.scala 19:72:@31855.4]
  assign _T_61891 = {storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7}; // @[Mux.scala 19:72:@31862.4]
  assign _T_61898 = {storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15}; // @[Mux.scala 19:72:@31869.4]
  assign _T_61899 = {storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,_T_61891}; // @[Mux.scala 19:72:@31870.4]
  assign _T_61901 = _T_2704 ? _T_61899 : 16'h0; // @[Mux.scala 19:72:@31871.4]
  assign _T_61916 = {storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,_T_61779}; // @[Mux.scala 19:72:@31886.4]
  assign _T_61918 = _T_2705 ? _T_61916 : 16'h0; // @[Mux.scala 19:72:@31887.4]
  assign _T_61933 = {storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,_T_61796}; // @[Mux.scala 19:72:@31902.4]
  assign _T_61935 = _T_2706 ? _T_61933 : 16'h0; // @[Mux.scala 19:72:@31903.4]
  assign _T_61950 = {storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,_T_61813}; // @[Mux.scala 19:72:@31918.4]
  assign _T_61952 = _T_2707 ? _T_61950 : 16'h0; // @[Mux.scala 19:72:@31919.4]
  assign _T_61967 = {storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,_T_61830}; // @[Mux.scala 19:72:@31934.4]
  assign _T_61969 = _T_2708 ? _T_61967 : 16'h0; // @[Mux.scala 19:72:@31935.4]
  assign _T_61984 = {storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,_T_61847}; // @[Mux.scala 19:72:@31950.4]
  assign _T_61986 = _T_2709 ? _T_61984 : 16'h0; // @[Mux.scala 19:72:@31951.4]
  assign _T_62001 = {storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,_T_61864}; // @[Mux.scala 19:72:@31966.4]
  assign _T_62003 = _T_2710 ? _T_62001 : 16'h0; // @[Mux.scala 19:72:@31967.4]
  assign _T_62018 = {storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,_T_61881}; // @[Mux.scala 19:72:@31982.4]
  assign _T_62020 = _T_2711 ? _T_62018 : 16'h0; // @[Mux.scala 19:72:@31983.4]
  assign _T_62035 = {storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,_T_61898}; // @[Mux.scala 19:72:@31998.4]
  assign _T_62037 = _T_2712 ? _T_62035 : 16'h0; // @[Mux.scala 19:72:@31999.4]
  assign _T_62038 = _T_61782 | _T_61799; // @[Mux.scala 19:72:@32000.4]
  assign _T_62039 = _T_62038 | _T_61816; // @[Mux.scala 19:72:@32001.4]
  assign _T_62040 = _T_62039 | _T_61833; // @[Mux.scala 19:72:@32002.4]
  assign _T_62041 = _T_62040 | _T_61850; // @[Mux.scala 19:72:@32003.4]
  assign _T_62042 = _T_62041 | _T_61867; // @[Mux.scala 19:72:@32004.4]
  assign _T_62043 = _T_62042 | _T_61884; // @[Mux.scala 19:72:@32005.4]
  assign _T_62044 = _T_62043 | _T_61901; // @[Mux.scala 19:72:@32006.4]
  assign _T_62045 = _T_62044 | _T_61918; // @[Mux.scala 19:72:@32007.4]
  assign _T_62046 = _T_62045 | _T_61935; // @[Mux.scala 19:72:@32008.4]
  assign _T_62047 = _T_62046 | _T_61952; // @[Mux.scala 19:72:@32009.4]
  assign _T_62048 = _T_62047 | _T_61969; // @[Mux.scala 19:72:@32010.4]
  assign _T_62049 = _T_62048 | _T_61986; // @[Mux.scala 19:72:@32011.4]
  assign _T_62050 = _T_62049 | _T_62003; // @[Mux.scala 19:72:@32012.4]
  assign _T_62051 = _T_62050 | _T_62020; // @[Mux.scala 19:72:@32013.4]
  assign _T_62052 = _T_62051 | _T_62037; // @[Mux.scala 19:72:@32014.4]
  assign _T_62630 = {storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0}; // @[Mux.scala 19:72:@32364.4]
  assign _T_62637 = {storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8}; // @[Mux.scala 19:72:@32371.4]
  assign _T_62638 = {storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,_T_62630}; // @[Mux.scala 19:72:@32372.4]
  assign _T_62640 = _T_2697 ? _T_62638 : 16'h0; // @[Mux.scala 19:72:@32373.4]
  assign _T_62647 = {storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1}; // @[Mux.scala 19:72:@32380.4]
  assign _T_62654 = {storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9}; // @[Mux.scala 19:72:@32387.4]
  assign _T_62655 = {storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,_T_62647}; // @[Mux.scala 19:72:@32388.4]
  assign _T_62657 = _T_2698 ? _T_62655 : 16'h0; // @[Mux.scala 19:72:@32389.4]
  assign _T_62664 = {storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2}; // @[Mux.scala 19:72:@32396.4]
  assign _T_62671 = {storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10}; // @[Mux.scala 19:72:@32403.4]
  assign _T_62672 = {storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,_T_62664}; // @[Mux.scala 19:72:@32404.4]
  assign _T_62674 = _T_2699 ? _T_62672 : 16'h0; // @[Mux.scala 19:72:@32405.4]
  assign _T_62681 = {storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3}; // @[Mux.scala 19:72:@32412.4]
  assign _T_62688 = {storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11}; // @[Mux.scala 19:72:@32419.4]
  assign _T_62689 = {storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,_T_62681}; // @[Mux.scala 19:72:@32420.4]
  assign _T_62691 = _T_2700 ? _T_62689 : 16'h0; // @[Mux.scala 19:72:@32421.4]
  assign _T_62698 = {storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4}; // @[Mux.scala 19:72:@32428.4]
  assign _T_62705 = {storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12}; // @[Mux.scala 19:72:@32435.4]
  assign _T_62706 = {storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,_T_62698}; // @[Mux.scala 19:72:@32436.4]
  assign _T_62708 = _T_2701 ? _T_62706 : 16'h0; // @[Mux.scala 19:72:@32437.4]
  assign _T_62715 = {storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5}; // @[Mux.scala 19:72:@32444.4]
  assign _T_62722 = {storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13}; // @[Mux.scala 19:72:@32451.4]
  assign _T_62723 = {storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,_T_62715}; // @[Mux.scala 19:72:@32452.4]
  assign _T_62725 = _T_2702 ? _T_62723 : 16'h0; // @[Mux.scala 19:72:@32453.4]
  assign _T_62732 = {storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6}; // @[Mux.scala 19:72:@32460.4]
  assign _T_62739 = {storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14}; // @[Mux.scala 19:72:@32467.4]
  assign _T_62740 = {storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,_T_62732}; // @[Mux.scala 19:72:@32468.4]
  assign _T_62742 = _T_2703 ? _T_62740 : 16'h0; // @[Mux.scala 19:72:@32469.4]
  assign _T_62749 = {storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7}; // @[Mux.scala 19:72:@32476.4]
  assign _T_62756 = {storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15}; // @[Mux.scala 19:72:@32483.4]
  assign _T_62757 = {storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,_T_62749}; // @[Mux.scala 19:72:@32484.4]
  assign _T_62759 = _T_2704 ? _T_62757 : 16'h0; // @[Mux.scala 19:72:@32485.4]
  assign _T_62774 = {storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,_T_62637}; // @[Mux.scala 19:72:@32500.4]
  assign _T_62776 = _T_2705 ? _T_62774 : 16'h0; // @[Mux.scala 19:72:@32501.4]
  assign _T_62791 = {storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,_T_62654}; // @[Mux.scala 19:72:@32516.4]
  assign _T_62793 = _T_2706 ? _T_62791 : 16'h0; // @[Mux.scala 19:72:@32517.4]
  assign _T_62808 = {storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,_T_62671}; // @[Mux.scala 19:72:@32532.4]
  assign _T_62810 = _T_2707 ? _T_62808 : 16'h0; // @[Mux.scala 19:72:@32533.4]
  assign _T_62825 = {storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,_T_62688}; // @[Mux.scala 19:72:@32548.4]
  assign _T_62827 = _T_2708 ? _T_62825 : 16'h0; // @[Mux.scala 19:72:@32549.4]
  assign _T_62842 = {storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,_T_62705}; // @[Mux.scala 19:72:@32564.4]
  assign _T_62844 = _T_2709 ? _T_62842 : 16'h0; // @[Mux.scala 19:72:@32565.4]
  assign _T_62859 = {storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,_T_62722}; // @[Mux.scala 19:72:@32580.4]
  assign _T_62861 = _T_2710 ? _T_62859 : 16'h0; // @[Mux.scala 19:72:@32581.4]
  assign _T_62876 = {storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,_T_62739}; // @[Mux.scala 19:72:@32596.4]
  assign _T_62878 = _T_2711 ? _T_62876 : 16'h0; // @[Mux.scala 19:72:@32597.4]
  assign _T_62893 = {storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,_T_62756}; // @[Mux.scala 19:72:@32612.4]
  assign _T_62895 = _T_2712 ? _T_62893 : 16'h0; // @[Mux.scala 19:72:@32613.4]
  assign _T_62896 = _T_62640 | _T_62657; // @[Mux.scala 19:72:@32614.4]
  assign _T_62897 = _T_62896 | _T_62674; // @[Mux.scala 19:72:@32615.4]
  assign _T_62898 = _T_62897 | _T_62691; // @[Mux.scala 19:72:@32616.4]
  assign _T_62899 = _T_62898 | _T_62708; // @[Mux.scala 19:72:@32617.4]
  assign _T_62900 = _T_62899 | _T_62725; // @[Mux.scala 19:72:@32618.4]
  assign _T_62901 = _T_62900 | _T_62742; // @[Mux.scala 19:72:@32619.4]
  assign _T_62902 = _T_62901 | _T_62759; // @[Mux.scala 19:72:@32620.4]
  assign _T_62903 = _T_62902 | _T_62776; // @[Mux.scala 19:72:@32621.4]
  assign _T_62904 = _T_62903 | _T_62793; // @[Mux.scala 19:72:@32622.4]
  assign _T_62905 = _T_62904 | _T_62810; // @[Mux.scala 19:72:@32623.4]
  assign _T_62906 = _T_62905 | _T_62827; // @[Mux.scala 19:72:@32624.4]
  assign _T_62907 = _T_62906 | _T_62844; // @[Mux.scala 19:72:@32625.4]
  assign _T_62908 = _T_62907 | _T_62861; // @[Mux.scala 19:72:@32626.4]
  assign _T_62909 = _T_62908 | _T_62878; // @[Mux.scala 19:72:@32627.4]
  assign _T_62910 = _T_62909 | _T_62895; // @[Mux.scala 19:72:@32628.4]
  assign _T_63488 = {storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0}; // @[Mux.scala 19:72:@32978.4]
  assign _T_63495 = {storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8}; // @[Mux.scala 19:72:@32985.4]
  assign _T_63496 = {storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,_T_63488}; // @[Mux.scala 19:72:@32986.4]
  assign _T_63498 = _T_2697 ? _T_63496 : 16'h0; // @[Mux.scala 19:72:@32987.4]
  assign _T_63505 = {storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1}; // @[Mux.scala 19:72:@32994.4]
  assign _T_63512 = {storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9}; // @[Mux.scala 19:72:@33001.4]
  assign _T_63513 = {storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,_T_63505}; // @[Mux.scala 19:72:@33002.4]
  assign _T_63515 = _T_2698 ? _T_63513 : 16'h0; // @[Mux.scala 19:72:@33003.4]
  assign _T_63522 = {storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2}; // @[Mux.scala 19:72:@33010.4]
  assign _T_63529 = {storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10}; // @[Mux.scala 19:72:@33017.4]
  assign _T_63530 = {storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,_T_63522}; // @[Mux.scala 19:72:@33018.4]
  assign _T_63532 = _T_2699 ? _T_63530 : 16'h0; // @[Mux.scala 19:72:@33019.4]
  assign _T_63539 = {storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3}; // @[Mux.scala 19:72:@33026.4]
  assign _T_63546 = {storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11}; // @[Mux.scala 19:72:@33033.4]
  assign _T_63547 = {storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,_T_63539}; // @[Mux.scala 19:72:@33034.4]
  assign _T_63549 = _T_2700 ? _T_63547 : 16'h0; // @[Mux.scala 19:72:@33035.4]
  assign _T_63556 = {storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4}; // @[Mux.scala 19:72:@33042.4]
  assign _T_63563 = {storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12}; // @[Mux.scala 19:72:@33049.4]
  assign _T_63564 = {storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,_T_63556}; // @[Mux.scala 19:72:@33050.4]
  assign _T_63566 = _T_2701 ? _T_63564 : 16'h0; // @[Mux.scala 19:72:@33051.4]
  assign _T_63573 = {storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5}; // @[Mux.scala 19:72:@33058.4]
  assign _T_63580 = {storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13}; // @[Mux.scala 19:72:@33065.4]
  assign _T_63581 = {storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,_T_63573}; // @[Mux.scala 19:72:@33066.4]
  assign _T_63583 = _T_2702 ? _T_63581 : 16'h0; // @[Mux.scala 19:72:@33067.4]
  assign _T_63590 = {storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6}; // @[Mux.scala 19:72:@33074.4]
  assign _T_63597 = {storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14}; // @[Mux.scala 19:72:@33081.4]
  assign _T_63598 = {storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,_T_63590}; // @[Mux.scala 19:72:@33082.4]
  assign _T_63600 = _T_2703 ? _T_63598 : 16'h0; // @[Mux.scala 19:72:@33083.4]
  assign _T_63607 = {storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7}; // @[Mux.scala 19:72:@33090.4]
  assign _T_63614 = {storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15}; // @[Mux.scala 19:72:@33097.4]
  assign _T_63615 = {storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,_T_63607}; // @[Mux.scala 19:72:@33098.4]
  assign _T_63617 = _T_2704 ? _T_63615 : 16'h0; // @[Mux.scala 19:72:@33099.4]
  assign _T_63632 = {storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,_T_63495}; // @[Mux.scala 19:72:@33114.4]
  assign _T_63634 = _T_2705 ? _T_63632 : 16'h0; // @[Mux.scala 19:72:@33115.4]
  assign _T_63649 = {storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,_T_63512}; // @[Mux.scala 19:72:@33130.4]
  assign _T_63651 = _T_2706 ? _T_63649 : 16'h0; // @[Mux.scala 19:72:@33131.4]
  assign _T_63666 = {storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,_T_63529}; // @[Mux.scala 19:72:@33146.4]
  assign _T_63668 = _T_2707 ? _T_63666 : 16'h0; // @[Mux.scala 19:72:@33147.4]
  assign _T_63683 = {storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,_T_63546}; // @[Mux.scala 19:72:@33162.4]
  assign _T_63685 = _T_2708 ? _T_63683 : 16'h0; // @[Mux.scala 19:72:@33163.4]
  assign _T_63700 = {storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,_T_63563}; // @[Mux.scala 19:72:@33178.4]
  assign _T_63702 = _T_2709 ? _T_63700 : 16'h0; // @[Mux.scala 19:72:@33179.4]
  assign _T_63717 = {storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,_T_63580}; // @[Mux.scala 19:72:@33194.4]
  assign _T_63719 = _T_2710 ? _T_63717 : 16'h0; // @[Mux.scala 19:72:@33195.4]
  assign _T_63734 = {storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,_T_63597}; // @[Mux.scala 19:72:@33210.4]
  assign _T_63736 = _T_2711 ? _T_63734 : 16'h0; // @[Mux.scala 19:72:@33211.4]
  assign _T_63751 = {storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,_T_63614}; // @[Mux.scala 19:72:@33226.4]
  assign _T_63753 = _T_2712 ? _T_63751 : 16'h0; // @[Mux.scala 19:72:@33227.4]
  assign _T_63754 = _T_63498 | _T_63515; // @[Mux.scala 19:72:@33228.4]
  assign _T_63755 = _T_63754 | _T_63532; // @[Mux.scala 19:72:@33229.4]
  assign _T_63756 = _T_63755 | _T_63549; // @[Mux.scala 19:72:@33230.4]
  assign _T_63757 = _T_63756 | _T_63566; // @[Mux.scala 19:72:@33231.4]
  assign _T_63758 = _T_63757 | _T_63583; // @[Mux.scala 19:72:@33232.4]
  assign _T_63759 = _T_63758 | _T_63600; // @[Mux.scala 19:72:@33233.4]
  assign _T_63760 = _T_63759 | _T_63617; // @[Mux.scala 19:72:@33234.4]
  assign _T_63761 = _T_63760 | _T_63634; // @[Mux.scala 19:72:@33235.4]
  assign _T_63762 = _T_63761 | _T_63651; // @[Mux.scala 19:72:@33236.4]
  assign _T_63763 = _T_63762 | _T_63668; // @[Mux.scala 19:72:@33237.4]
  assign _T_63764 = _T_63763 | _T_63685; // @[Mux.scala 19:72:@33238.4]
  assign _T_63765 = _T_63764 | _T_63702; // @[Mux.scala 19:72:@33239.4]
  assign _T_63766 = _T_63765 | _T_63719; // @[Mux.scala 19:72:@33240.4]
  assign _T_63767 = _T_63766 | _T_63736; // @[Mux.scala 19:72:@33241.4]
  assign _T_63768 = _T_63767 | _T_63753; // @[Mux.scala 19:72:@33242.4]
  assign _T_64346 = {storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0}; // @[Mux.scala 19:72:@33592.4]
  assign _T_64353 = {storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8}; // @[Mux.scala 19:72:@33599.4]
  assign _T_64354 = {storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,_T_64346}; // @[Mux.scala 19:72:@33600.4]
  assign _T_64356 = _T_2697 ? _T_64354 : 16'h0; // @[Mux.scala 19:72:@33601.4]
  assign _T_64363 = {storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1}; // @[Mux.scala 19:72:@33608.4]
  assign _T_64370 = {storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9}; // @[Mux.scala 19:72:@33615.4]
  assign _T_64371 = {storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,_T_64363}; // @[Mux.scala 19:72:@33616.4]
  assign _T_64373 = _T_2698 ? _T_64371 : 16'h0; // @[Mux.scala 19:72:@33617.4]
  assign _T_64380 = {storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2}; // @[Mux.scala 19:72:@33624.4]
  assign _T_64387 = {storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10}; // @[Mux.scala 19:72:@33631.4]
  assign _T_64388 = {storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,_T_64380}; // @[Mux.scala 19:72:@33632.4]
  assign _T_64390 = _T_2699 ? _T_64388 : 16'h0; // @[Mux.scala 19:72:@33633.4]
  assign _T_64397 = {storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3}; // @[Mux.scala 19:72:@33640.4]
  assign _T_64404 = {storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11}; // @[Mux.scala 19:72:@33647.4]
  assign _T_64405 = {storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,_T_64397}; // @[Mux.scala 19:72:@33648.4]
  assign _T_64407 = _T_2700 ? _T_64405 : 16'h0; // @[Mux.scala 19:72:@33649.4]
  assign _T_64414 = {storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4}; // @[Mux.scala 19:72:@33656.4]
  assign _T_64421 = {storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12}; // @[Mux.scala 19:72:@33663.4]
  assign _T_64422 = {storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,_T_64414}; // @[Mux.scala 19:72:@33664.4]
  assign _T_64424 = _T_2701 ? _T_64422 : 16'h0; // @[Mux.scala 19:72:@33665.4]
  assign _T_64431 = {storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5}; // @[Mux.scala 19:72:@33672.4]
  assign _T_64438 = {storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13}; // @[Mux.scala 19:72:@33679.4]
  assign _T_64439 = {storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,_T_64431}; // @[Mux.scala 19:72:@33680.4]
  assign _T_64441 = _T_2702 ? _T_64439 : 16'h0; // @[Mux.scala 19:72:@33681.4]
  assign _T_64448 = {storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6}; // @[Mux.scala 19:72:@33688.4]
  assign _T_64455 = {storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14}; // @[Mux.scala 19:72:@33695.4]
  assign _T_64456 = {storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,_T_64448}; // @[Mux.scala 19:72:@33696.4]
  assign _T_64458 = _T_2703 ? _T_64456 : 16'h0; // @[Mux.scala 19:72:@33697.4]
  assign _T_64465 = {storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7}; // @[Mux.scala 19:72:@33704.4]
  assign _T_64472 = {storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15}; // @[Mux.scala 19:72:@33711.4]
  assign _T_64473 = {storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,_T_64465}; // @[Mux.scala 19:72:@33712.4]
  assign _T_64475 = _T_2704 ? _T_64473 : 16'h0; // @[Mux.scala 19:72:@33713.4]
  assign _T_64490 = {storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,_T_64353}; // @[Mux.scala 19:72:@33728.4]
  assign _T_64492 = _T_2705 ? _T_64490 : 16'h0; // @[Mux.scala 19:72:@33729.4]
  assign _T_64507 = {storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,_T_64370}; // @[Mux.scala 19:72:@33744.4]
  assign _T_64509 = _T_2706 ? _T_64507 : 16'h0; // @[Mux.scala 19:72:@33745.4]
  assign _T_64524 = {storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,_T_64387}; // @[Mux.scala 19:72:@33760.4]
  assign _T_64526 = _T_2707 ? _T_64524 : 16'h0; // @[Mux.scala 19:72:@33761.4]
  assign _T_64541 = {storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,_T_64404}; // @[Mux.scala 19:72:@33776.4]
  assign _T_64543 = _T_2708 ? _T_64541 : 16'h0; // @[Mux.scala 19:72:@33777.4]
  assign _T_64558 = {storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,_T_64421}; // @[Mux.scala 19:72:@33792.4]
  assign _T_64560 = _T_2709 ? _T_64558 : 16'h0; // @[Mux.scala 19:72:@33793.4]
  assign _T_64575 = {storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,_T_64438}; // @[Mux.scala 19:72:@33808.4]
  assign _T_64577 = _T_2710 ? _T_64575 : 16'h0; // @[Mux.scala 19:72:@33809.4]
  assign _T_64592 = {storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,_T_64455}; // @[Mux.scala 19:72:@33824.4]
  assign _T_64594 = _T_2711 ? _T_64592 : 16'h0; // @[Mux.scala 19:72:@33825.4]
  assign _T_64609 = {storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,_T_64472}; // @[Mux.scala 19:72:@33840.4]
  assign _T_64611 = _T_2712 ? _T_64609 : 16'h0; // @[Mux.scala 19:72:@33841.4]
  assign _T_64612 = _T_64356 | _T_64373; // @[Mux.scala 19:72:@33842.4]
  assign _T_64613 = _T_64612 | _T_64390; // @[Mux.scala 19:72:@33843.4]
  assign _T_64614 = _T_64613 | _T_64407; // @[Mux.scala 19:72:@33844.4]
  assign _T_64615 = _T_64614 | _T_64424; // @[Mux.scala 19:72:@33845.4]
  assign _T_64616 = _T_64615 | _T_64441; // @[Mux.scala 19:72:@33846.4]
  assign _T_64617 = _T_64616 | _T_64458; // @[Mux.scala 19:72:@33847.4]
  assign _T_64618 = _T_64617 | _T_64475; // @[Mux.scala 19:72:@33848.4]
  assign _T_64619 = _T_64618 | _T_64492; // @[Mux.scala 19:72:@33849.4]
  assign _T_64620 = _T_64619 | _T_64509; // @[Mux.scala 19:72:@33850.4]
  assign _T_64621 = _T_64620 | _T_64526; // @[Mux.scala 19:72:@33851.4]
  assign _T_64622 = _T_64621 | _T_64543; // @[Mux.scala 19:72:@33852.4]
  assign _T_64623 = _T_64622 | _T_64560; // @[Mux.scala 19:72:@33853.4]
  assign _T_64624 = _T_64623 | _T_64577; // @[Mux.scala 19:72:@33854.4]
  assign _T_64625 = _T_64624 | _T_64594; // @[Mux.scala 19:72:@33855.4]
  assign _T_64626 = _T_64625 | _T_64611; // @[Mux.scala 19:72:@33856.4]
  assign _T_65204 = {storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0}; // @[Mux.scala 19:72:@34206.4]
  assign _T_65211 = {storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8}; // @[Mux.scala 19:72:@34213.4]
  assign _T_65212 = {storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,_T_65204}; // @[Mux.scala 19:72:@34214.4]
  assign _T_65214 = _T_2697 ? _T_65212 : 16'h0; // @[Mux.scala 19:72:@34215.4]
  assign _T_65221 = {storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1}; // @[Mux.scala 19:72:@34222.4]
  assign _T_65228 = {storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9}; // @[Mux.scala 19:72:@34229.4]
  assign _T_65229 = {storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,_T_65221}; // @[Mux.scala 19:72:@34230.4]
  assign _T_65231 = _T_2698 ? _T_65229 : 16'h0; // @[Mux.scala 19:72:@34231.4]
  assign _T_65238 = {storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2}; // @[Mux.scala 19:72:@34238.4]
  assign _T_65245 = {storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10}; // @[Mux.scala 19:72:@34245.4]
  assign _T_65246 = {storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,_T_65238}; // @[Mux.scala 19:72:@34246.4]
  assign _T_65248 = _T_2699 ? _T_65246 : 16'h0; // @[Mux.scala 19:72:@34247.4]
  assign _T_65255 = {storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3}; // @[Mux.scala 19:72:@34254.4]
  assign _T_65262 = {storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11}; // @[Mux.scala 19:72:@34261.4]
  assign _T_65263 = {storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,_T_65255}; // @[Mux.scala 19:72:@34262.4]
  assign _T_65265 = _T_2700 ? _T_65263 : 16'h0; // @[Mux.scala 19:72:@34263.4]
  assign _T_65272 = {storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4}; // @[Mux.scala 19:72:@34270.4]
  assign _T_65279 = {storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12}; // @[Mux.scala 19:72:@34277.4]
  assign _T_65280 = {storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,_T_65272}; // @[Mux.scala 19:72:@34278.4]
  assign _T_65282 = _T_2701 ? _T_65280 : 16'h0; // @[Mux.scala 19:72:@34279.4]
  assign _T_65289 = {storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5}; // @[Mux.scala 19:72:@34286.4]
  assign _T_65296 = {storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13}; // @[Mux.scala 19:72:@34293.4]
  assign _T_65297 = {storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,_T_65289}; // @[Mux.scala 19:72:@34294.4]
  assign _T_65299 = _T_2702 ? _T_65297 : 16'h0; // @[Mux.scala 19:72:@34295.4]
  assign _T_65306 = {storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6}; // @[Mux.scala 19:72:@34302.4]
  assign _T_65313 = {storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14}; // @[Mux.scala 19:72:@34309.4]
  assign _T_65314 = {storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,_T_65306}; // @[Mux.scala 19:72:@34310.4]
  assign _T_65316 = _T_2703 ? _T_65314 : 16'h0; // @[Mux.scala 19:72:@34311.4]
  assign _T_65323 = {storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7}; // @[Mux.scala 19:72:@34318.4]
  assign _T_65330 = {storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15}; // @[Mux.scala 19:72:@34325.4]
  assign _T_65331 = {storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,_T_65323}; // @[Mux.scala 19:72:@34326.4]
  assign _T_65333 = _T_2704 ? _T_65331 : 16'h0; // @[Mux.scala 19:72:@34327.4]
  assign _T_65348 = {storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,_T_65211}; // @[Mux.scala 19:72:@34342.4]
  assign _T_65350 = _T_2705 ? _T_65348 : 16'h0; // @[Mux.scala 19:72:@34343.4]
  assign _T_65365 = {storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,_T_65228}; // @[Mux.scala 19:72:@34358.4]
  assign _T_65367 = _T_2706 ? _T_65365 : 16'h0; // @[Mux.scala 19:72:@34359.4]
  assign _T_65382 = {storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,_T_65245}; // @[Mux.scala 19:72:@34374.4]
  assign _T_65384 = _T_2707 ? _T_65382 : 16'h0; // @[Mux.scala 19:72:@34375.4]
  assign _T_65399 = {storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,_T_65262}; // @[Mux.scala 19:72:@34390.4]
  assign _T_65401 = _T_2708 ? _T_65399 : 16'h0; // @[Mux.scala 19:72:@34391.4]
  assign _T_65416 = {storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,_T_65279}; // @[Mux.scala 19:72:@34406.4]
  assign _T_65418 = _T_2709 ? _T_65416 : 16'h0; // @[Mux.scala 19:72:@34407.4]
  assign _T_65433 = {storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,_T_65296}; // @[Mux.scala 19:72:@34422.4]
  assign _T_65435 = _T_2710 ? _T_65433 : 16'h0; // @[Mux.scala 19:72:@34423.4]
  assign _T_65450 = {storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,_T_65313}; // @[Mux.scala 19:72:@34438.4]
  assign _T_65452 = _T_2711 ? _T_65450 : 16'h0; // @[Mux.scala 19:72:@34439.4]
  assign _T_65467 = {storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,_T_65330}; // @[Mux.scala 19:72:@34454.4]
  assign _T_65469 = _T_2712 ? _T_65467 : 16'h0; // @[Mux.scala 19:72:@34455.4]
  assign _T_65470 = _T_65214 | _T_65231; // @[Mux.scala 19:72:@34456.4]
  assign _T_65471 = _T_65470 | _T_65248; // @[Mux.scala 19:72:@34457.4]
  assign _T_65472 = _T_65471 | _T_65265; // @[Mux.scala 19:72:@34458.4]
  assign _T_65473 = _T_65472 | _T_65282; // @[Mux.scala 19:72:@34459.4]
  assign _T_65474 = _T_65473 | _T_65299; // @[Mux.scala 19:72:@34460.4]
  assign _T_65475 = _T_65474 | _T_65316; // @[Mux.scala 19:72:@34461.4]
  assign _T_65476 = _T_65475 | _T_65333; // @[Mux.scala 19:72:@34462.4]
  assign _T_65477 = _T_65476 | _T_65350; // @[Mux.scala 19:72:@34463.4]
  assign _T_65478 = _T_65477 | _T_65367; // @[Mux.scala 19:72:@34464.4]
  assign _T_65479 = _T_65478 | _T_65384; // @[Mux.scala 19:72:@34465.4]
  assign _T_65480 = _T_65479 | _T_65401; // @[Mux.scala 19:72:@34466.4]
  assign _T_65481 = _T_65480 | _T_65418; // @[Mux.scala 19:72:@34467.4]
  assign _T_65482 = _T_65481 | _T_65435; // @[Mux.scala 19:72:@34468.4]
  assign _T_65483 = _T_65482 | _T_65452; // @[Mux.scala 19:72:@34469.4]
  assign _T_65484 = _T_65483 | _T_65469; // @[Mux.scala 19:72:@34470.4]
  assign _T_88276 = conflictPReg_0_2 ? 2'h2 : {{1'd0}, conflictPReg_0_1}; // @[LoadQueue.scala 191:60:@35143.4]
  assign _T_88277 = conflictPReg_0_3 ? 2'h3 : _T_88276; // @[LoadQueue.scala 191:60:@35144.4]
  assign _T_88278 = conflictPReg_0_4 ? 3'h4 : {{1'd0}, _T_88277}; // @[LoadQueue.scala 191:60:@35145.4]
  assign _T_88279 = conflictPReg_0_5 ? 3'h5 : _T_88278; // @[LoadQueue.scala 191:60:@35146.4]
  assign _T_88280 = conflictPReg_0_6 ? 3'h6 : _T_88279; // @[LoadQueue.scala 191:60:@35147.4]
  assign _T_88281 = conflictPReg_0_7 ? 3'h7 : _T_88280; // @[LoadQueue.scala 191:60:@35148.4]
  assign _T_88282 = conflictPReg_0_8 ? 4'h8 : {{1'd0}, _T_88281}; // @[LoadQueue.scala 191:60:@35149.4]
  assign _T_88283 = conflictPReg_0_9 ? 4'h9 : _T_88282; // @[LoadQueue.scala 191:60:@35150.4]
  assign _T_88284 = conflictPReg_0_10 ? 4'ha : _T_88283; // @[LoadQueue.scala 191:60:@35151.4]
  assign _T_88285 = conflictPReg_0_11 ? 4'hb : _T_88284; // @[LoadQueue.scala 191:60:@35152.4]
  assign _T_88286 = conflictPReg_0_12 ? 4'hc : _T_88285; // @[LoadQueue.scala 191:60:@35153.4]
  assign _T_88287 = conflictPReg_0_13 ? 4'hd : _T_88286; // @[LoadQueue.scala 191:60:@35154.4]
  assign _T_88288 = conflictPReg_0_14 ? 4'he : _T_88287; // @[LoadQueue.scala 191:60:@35155.4]
  assign _T_88289 = conflictPReg_0_15 ? 4'hf : _T_88288; // @[LoadQueue.scala 191:60:@35156.4]
  assign _T_88292 = conflictPReg_0_0 | conflictPReg_0_1; // @[LoadQueue.scala 192:43:@35158.4]
  assign _T_88293 = _T_88292 | conflictPReg_0_2; // @[LoadQueue.scala 192:43:@35159.4]
  assign _T_88294 = _T_88293 | conflictPReg_0_3; // @[LoadQueue.scala 192:43:@35160.4]
  assign _T_88295 = _T_88294 | conflictPReg_0_4; // @[LoadQueue.scala 192:43:@35161.4]
  assign _T_88296 = _T_88295 | conflictPReg_0_5; // @[LoadQueue.scala 192:43:@35162.4]
  assign _T_88297 = _T_88296 | conflictPReg_0_6; // @[LoadQueue.scala 192:43:@35163.4]
  assign _T_88298 = _T_88297 | conflictPReg_0_7; // @[LoadQueue.scala 192:43:@35164.4]
  assign _T_88299 = _T_88298 | conflictPReg_0_8; // @[LoadQueue.scala 192:43:@35165.4]
  assign _T_88300 = _T_88299 | conflictPReg_0_9; // @[LoadQueue.scala 192:43:@35166.4]
  assign _T_88301 = _T_88300 | conflictPReg_0_10; // @[LoadQueue.scala 192:43:@35167.4]
  assign _T_88302 = _T_88301 | conflictPReg_0_11; // @[LoadQueue.scala 192:43:@35168.4]
  assign _T_88303 = _T_88302 | conflictPReg_0_12; // @[LoadQueue.scala 192:43:@35169.4]
  assign _T_88304 = _T_88303 | conflictPReg_0_13; // @[LoadQueue.scala 192:43:@35170.4]
  assign _T_88305 = _T_88304 | conflictPReg_0_14; // @[LoadQueue.scala 192:43:@35171.4]
  assign _T_88306 = _T_88305 | conflictPReg_0_15; // @[LoadQueue.scala 192:43:@35172.4]
  assign _GEN_864 = 4'h0 == _T_88289; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_865 = 4'h1 == _T_88289; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_866 = 4'h2 == _T_88289; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_867 = 4'h3 == _T_88289; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_868 = 4'h4 == _T_88289; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_869 = 4'h5 == _T_88289; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_870 = 4'h6 == _T_88289; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_871 = 4'h7 == _T_88289; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_872 = 4'h8 == _T_88289; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_873 = 4'h9 == _T_88289; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_874 = 4'ha == _T_88289; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_875 = 4'hb == _T_88289; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_876 = 4'hc == _T_88289; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_877 = 4'hd == _T_88289; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_878 = 4'he == _T_88289; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_879 = 4'hf == _T_88289; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_881 = 4'h1 == _T_88289 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_882 = 4'h2 == _T_88289 ? shiftedStoreDataKnownPReg_2 : _GEN_881; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_883 = 4'h3 == _T_88289 ? shiftedStoreDataKnownPReg_3 : _GEN_882; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_884 = 4'h4 == _T_88289 ? shiftedStoreDataKnownPReg_4 : _GEN_883; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_885 = 4'h5 == _T_88289 ? shiftedStoreDataKnownPReg_5 : _GEN_884; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_886 = 4'h6 == _T_88289 ? shiftedStoreDataKnownPReg_6 : _GEN_885; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_887 = 4'h7 == _T_88289 ? shiftedStoreDataKnownPReg_7 : _GEN_886; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_888 = 4'h8 == _T_88289 ? shiftedStoreDataKnownPReg_8 : _GEN_887; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_889 = 4'h9 == _T_88289 ? shiftedStoreDataKnownPReg_9 : _GEN_888; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_890 = 4'ha == _T_88289 ? shiftedStoreDataKnownPReg_10 : _GEN_889; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_891 = 4'hb == _T_88289 ? shiftedStoreDataKnownPReg_11 : _GEN_890; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_892 = 4'hc == _T_88289 ? shiftedStoreDataKnownPReg_12 : _GEN_891; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_893 = 4'hd == _T_88289 ? shiftedStoreDataKnownPReg_13 : _GEN_892; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_894 = 4'he == _T_88289 ? shiftedStoreDataKnownPReg_14 : _GEN_893; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_895 = 4'hf == _T_88289 ? shiftedStoreDataKnownPReg_15 : _GEN_894; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_897 = 4'h1 == _T_88289 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_898 = 4'h2 == _T_88289 ? shiftedStoreDataQPreg_2 : _GEN_897; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_899 = 4'h3 == _T_88289 ? shiftedStoreDataQPreg_3 : _GEN_898; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_900 = 4'h4 == _T_88289 ? shiftedStoreDataQPreg_4 : _GEN_899; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_901 = 4'h5 == _T_88289 ? shiftedStoreDataQPreg_5 : _GEN_900; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_902 = 4'h6 == _T_88289 ? shiftedStoreDataQPreg_6 : _GEN_901; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_903 = 4'h7 == _T_88289 ? shiftedStoreDataQPreg_7 : _GEN_902; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_904 = 4'h8 == _T_88289 ? shiftedStoreDataQPreg_8 : _GEN_903; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_905 = 4'h9 == _T_88289 ? shiftedStoreDataQPreg_9 : _GEN_904; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_906 = 4'ha == _T_88289 ? shiftedStoreDataQPreg_10 : _GEN_905; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_907 = 4'hb == _T_88289 ? shiftedStoreDataQPreg_11 : _GEN_906; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_908 = 4'hc == _T_88289 ? shiftedStoreDataQPreg_12 : _GEN_907; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_909 = 4'hd == _T_88289 ? shiftedStoreDataQPreg_13 : _GEN_908; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_910 = 4'he == _T_88289 ? shiftedStoreDataQPreg_14 : _GEN_909; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_911 = 4'hf == _T_88289 ? shiftedStoreDataQPreg_15 : _GEN_910; // @[LoadQueue.scala 195:31:@35176.6]
  assign lastConflict_0_0 = _T_88306 ? _GEN_864 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_1 = _T_88306 ? _GEN_865 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_2 = _T_88306 ? _GEN_866 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_3 = _T_88306 ? _GEN_867 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_4 = _T_88306 ? _GEN_868 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_5 = _T_88306 ? _GEN_869 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_6 = _T_88306 ? _GEN_870 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_7 = _T_88306 ? _GEN_871 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_8 = _T_88306 ? _GEN_872 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_9 = _T_88306 ? _GEN_873 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_10 = _T_88306 ? _GEN_874 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_11 = _T_88306 ? _GEN_875 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_12 = _T_88306 ? _GEN_876 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_13 = _T_88306 ? _GEN_877 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_14 = _T_88306 ? _GEN_878 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_15 = _T_88306 ? _GEN_879 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign canBypass_0 = _T_88306 ? _GEN_895 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign bypassVal_0 = _T_88306 ? _GEN_911 : 32'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign _T_88412 = conflictPReg_1_2 ? 2'h2 : {{1'd0}, conflictPReg_1_1}; // @[LoadQueue.scala 191:60:@35230.4]
  assign _T_88413 = conflictPReg_1_3 ? 2'h3 : _T_88412; // @[LoadQueue.scala 191:60:@35231.4]
  assign _T_88414 = conflictPReg_1_4 ? 3'h4 : {{1'd0}, _T_88413}; // @[LoadQueue.scala 191:60:@35232.4]
  assign _T_88415 = conflictPReg_1_5 ? 3'h5 : _T_88414; // @[LoadQueue.scala 191:60:@35233.4]
  assign _T_88416 = conflictPReg_1_6 ? 3'h6 : _T_88415; // @[LoadQueue.scala 191:60:@35234.4]
  assign _T_88417 = conflictPReg_1_7 ? 3'h7 : _T_88416; // @[LoadQueue.scala 191:60:@35235.4]
  assign _T_88418 = conflictPReg_1_8 ? 4'h8 : {{1'd0}, _T_88417}; // @[LoadQueue.scala 191:60:@35236.4]
  assign _T_88419 = conflictPReg_1_9 ? 4'h9 : _T_88418; // @[LoadQueue.scala 191:60:@35237.4]
  assign _T_88420 = conflictPReg_1_10 ? 4'ha : _T_88419; // @[LoadQueue.scala 191:60:@35238.4]
  assign _T_88421 = conflictPReg_1_11 ? 4'hb : _T_88420; // @[LoadQueue.scala 191:60:@35239.4]
  assign _T_88422 = conflictPReg_1_12 ? 4'hc : _T_88421; // @[LoadQueue.scala 191:60:@35240.4]
  assign _T_88423 = conflictPReg_1_13 ? 4'hd : _T_88422; // @[LoadQueue.scala 191:60:@35241.4]
  assign _T_88424 = conflictPReg_1_14 ? 4'he : _T_88423; // @[LoadQueue.scala 191:60:@35242.4]
  assign _T_88425 = conflictPReg_1_15 ? 4'hf : _T_88424; // @[LoadQueue.scala 191:60:@35243.4]
  assign _T_88428 = conflictPReg_1_0 | conflictPReg_1_1; // @[LoadQueue.scala 192:43:@35245.4]
  assign _T_88429 = _T_88428 | conflictPReg_1_2; // @[LoadQueue.scala 192:43:@35246.4]
  assign _T_88430 = _T_88429 | conflictPReg_1_3; // @[LoadQueue.scala 192:43:@35247.4]
  assign _T_88431 = _T_88430 | conflictPReg_1_4; // @[LoadQueue.scala 192:43:@35248.4]
  assign _T_88432 = _T_88431 | conflictPReg_1_5; // @[LoadQueue.scala 192:43:@35249.4]
  assign _T_88433 = _T_88432 | conflictPReg_1_6; // @[LoadQueue.scala 192:43:@35250.4]
  assign _T_88434 = _T_88433 | conflictPReg_1_7; // @[LoadQueue.scala 192:43:@35251.4]
  assign _T_88435 = _T_88434 | conflictPReg_1_8; // @[LoadQueue.scala 192:43:@35252.4]
  assign _T_88436 = _T_88435 | conflictPReg_1_9; // @[LoadQueue.scala 192:43:@35253.4]
  assign _T_88437 = _T_88436 | conflictPReg_1_10; // @[LoadQueue.scala 192:43:@35254.4]
  assign _T_88438 = _T_88437 | conflictPReg_1_11; // @[LoadQueue.scala 192:43:@35255.4]
  assign _T_88439 = _T_88438 | conflictPReg_1_12; // @[LoadQueue.scala 192:43:@35256.4]
  assign _T_88440 = _T_88439 | conflictPReg_1_13; // @[LoadQueue.scala 192:43:@35257.4]
  assign _T_88441 = _T_88440 | conflictPReg_1_14; // @[LoadQueue.scala 192:43:@35258.4]
  assign _T_88442 = _T_88441 | conflictPReg_1_15; // @[LoadQueue.scala 192:43:@35259.4]
  assign _GEN_930 = 4'h0 == _T_88425; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_931 = 4'h1 == _T_88425; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_932 = 4'h2 == _T_88425; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_933 = 4'h3 == _T_88425; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_934 = 4'h4 == _T_88425; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_935 = 4'h5 == _T_88425; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_936 = 4'h6 == _T_88425; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_937 = 4'h7 == _T_88425; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_938 = 4'h8 == _T_88425; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_939 = 4'h9 == _T_88425; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_940 = 4'ha == _T_88425; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_941 = 4'hb == _T_88425; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_942 = 4'hc == _T_88425; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_943 = 4'hd == _T_88425; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_944 = 4'he == _T_88425; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_945 = 4'hf == _T_88425; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_947 = 4'h1 == _T_88425 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_948 = 4'h2 == _T_88425 ? shiftedStoreDataKnownPReg_2 : _GEN_947; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_949 = 4'h3 == _T_88425 ? shiftedStoreDataKnownPReg_3 : _GEN_948; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_950 = 4'h4 == _T_88425 ? shiftedStoreDataKnownPReg_4 : _GEN_949; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_951 = 4'h5 == _T_88425 ? shiftedStoreDataKnownPReg_5 : _GEN_950; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_952 = 4'h6 == _T_88425 ? shiftedStoreDataKnownPReg_6 : _GEN_951; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_953 = 4'h7 == _T_88425 ? shiftedStoreDataKnownPReg_7 : _GEN_952; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_954 = 4'h8 == _T_88425 ? shiftedStoreDataKnownPReg_8 : _GEN_953; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_955 = 4'h9 == _T_88425 ? shiftedStoreDataKnownPReg_9 : _GEN_954; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_956 = 4'ha == _T_88425 ? shiftedStoreDataKnownPReg_10 : _GEN_955; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_957 = 4'hb == _T_88425 ? shiftedStoreDataKnownPReg_11 : _GEN_956; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_958 = 4'hc == _T_88425 ? shiftedStoreDataKnownPReg_12 : _GEN_957; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_959 = 4'hd == _T_88425 ? shiftedStoreDataKnownPReg_13 : _GEN_958; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_960 = 4'he == _T_88425 ? shiftedStoreDataKnownPReg_14 : _GEN_959; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_961 = 4'hf == _T_88425 ? shiftedStoreDataKnownPReg_15 : _GEN_960; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_963 = 4'h1 == _T_88425 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_964 = 4'h2 == _T_88425 ? shiftedStoreDataQPreg_2 : _GEN_963; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_965 = 4'h3 == _T_88425 ? shiftedStoreDataQPreg_3 : _GEN_964; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_966 = 4'h4 == _T_88425 ? shiftedStoreDataQPreg_4 : _GEN_965; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_967 = 4'h5 == _T_88425 ? shiftedStoreDataQPreg_5 : _GEN_966; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_968 = 4'h6 == _T_88425 ? shiftedStoreDataQPreg_6 : _GEN_967; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_969 = 4'h7 == _T_88425 ? shiftedStoreDataQPreg_7 : _GEN_968; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_970 = 4'h8 == _T_88425 ? shiftedStoreDataQPreg_8 : _GEN_969; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_971 = 4'h9 == _T_88425 ? shiftedStoreDataQPreg_9 : _GEN_970; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_972 = 4'ha == _T_88425 ? shiftedStoreDataQPreg_10 : _GEN_971; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_973 = 4'hb == _T_88425 ? shiftedStoreDataQPreg_11 : _GEN_972; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_974 = 4'hc == _T_88425 ? shiftedStoreDataQPreg_12 : _GEN_973; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_975 = 4'hd == _T_88425 ? shiftedStoreDataQPreg_13 : _GEN_974; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_976 = 4'he == _T_88425 ? shiftedStoreDataQPreg_14 : _GEN_975; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_977 = 4'hf == _T_88425 ? shiftedStoreDataQPreg_15 : _GEN_976; // @[LoadQueue.scala 195:31:@35263.6]
  assign lastConflict_1_0 = _T_88442 ? _GEN_930 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_1 = _T_88442 ? _GEN_931 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_2 = _T_88442 ? _GEN_932 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_3 = _T_88442 ? _GEN_933 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_4 = _T_88442 ? _GEN_934 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_5 = _T_88442 ? _GEN_935 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_6 = _T_88442 ? _GEN_936 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_7 = _T_88442 ? _GEN_937 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_8 = _T_88442 ? _GEN_938 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_9 = _T_88442 ? _GEN_939 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_10 = _T_88442 ? _GEN_940 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_11 = _T_88442 ? _GEN_941 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_12 = _T_88442 ? _GEN_942 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_13 = _T_88442 ? _GEN_943 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_14 = _T_88442 ? _GEN_944 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_15 = _T_88442 ? _GEN_945 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign canBypass_1 = _T_88442 ? _GEN_961 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign bypassVal_1 = _T_88442 ? _GEN_977 : 32'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign _T_88548 = conflictPReg_2_2 ? 2'h2 : {{1'd0}, conflictPReg_2_1}; // @[LoadQueue.scala 191:60:@35317.4]
  assign _T_88549 = conflictPReg_2_3 ? 2'h3 : _T_88548; // @[LoadQueue.scala 191:60:@35318.4]
  assign _T_88550 = conflictPReg_2_4 ? 3'h4 : {{1'd0}, _T_88549}; // @[LoadQueue.scala 191:60:@35319.4]
  assign _T_88551 = conflictPReg_2_5 ? 3'h5 : _T_88550; // @[LoadQueue.scala 191:60:@35320.4]
  assign _T_88552 = conflictPReg_2_6 ? 3'h6 : _T_88551; // @[LoadQueue.scala 191:60:@35321.4]
  assign _T_88553 = conflictPReg_2_7 ? 3'h7 : _T_88552; // @[LoadQueue.scala 191:60:@35322.4]
  assign _T_88554 = conflictPReg_2_8 ? 4'h8 : {{1'd0}, _T_88553}; // @[LoadQueue.scala 191:60:@35323.4]
  assign _T_88555 = conflictPReg_2_9 ? 4'h9 : _T_88554; // @[LoadQueue.scala 191:60:@35324.4]
  assign _T_88556 = conflictPReg_2_10 ? 4'ha : _T_88555; // @[LoadQueue.scala 191:60:@35325.4]
  assign _T_88557 = conflictPReg_2_11 ? 4'hb : _T_88556; // @[LoadQueue.scala 191:60:@35326.4]
  assign _T_88558 = conflictPReg_2_12 ? 4'hc : _T_88557; // @[LoadQueue.scala 191:60:@35327.4]
  assign _T_88559 = conflictPReg_2_13 ? 4'hd : _T_88558; // @[LoadQueue.scala 191:60:@35328.4]
  assign _T_88560 = conflictPReg_2_14 ? 4'he : _T_88559; // @[LoadQueue.scala 191:60:@35329.4]
  assign _T_88561 = conflictPReg_2_15 ? 4'hf : _T_88560; // @[LoadQueue.scala 191:60:@35330.4]
  assign _T_88564 = conflictPReg_2_0 | conflictPReg_2_1; // @[LoadQueue.scala 192:43:@35332.4]
  assign _T_88565 = _T_88564 | conflictPReg_2_2; // @[LoadQueue.scala 192:43:@35333.4]
  assign _T_88566 = _T_88565 | conflictPReg_2_3; // @[LoadQueue.scala 192:43:@35334.4]
  assign _T_88567 = _T_88566 | conflictPReg_2_4; // @[LoadQueue.scala 192:43:@35335.4]
  assign _T_88568 = _T_88567 | conflictPReg_2_5; // @[LoadQueue.scala 192:43:@35336.4]
  assign _T_88569 = _T_88568 | conflictPReg_2_6; // @[LoadQueue.scala 192:43:@35337.4]
  assign _T_88570 = _T_88569 | conflictPReg_2_7; // @[LoadQueue.scala 192:43:@35338.4]
  assign _T_88571 = _T_88570 | conflictPReg_2_8; // @[LoadQueue.scala 192:43:@35339.4]
  assign _T_88572 = _T_88571 | conflictPReg_2_9; // @[LoadQueue.scala 192:43:@35340.4]
  assign _T_88573 = _T_88572 | conflictPReg_2_10; // @[LoadQueue.scala 192:43:@35341.4]
  assign _T_88574 = _T_88573 | conflictPReg_2_11; // @[LoadQueue.scala 192:43:@35342.4]
  assign _T_88575 = _T_88574 | conflictPReg_2_12; // @[LoadQueue.scala 192:43:@35343.4]
  assign _T_88576 = _T_88575 | conflictPReg_2_13; // @[LoadQueue.scala 192:43:@35344.4]
  assign _T_88577 = _T_88576 | conflictPReg_2_14; // @[LoadQueue.scala 192:43:@35345.4]
  assign _T_88578 = _T_88577 | conflictPReg_2_15; // @[LoadQueue.scala 192:43:@35346.4]
  assign _GEN_996 = 4'h0 == _T_88561; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_997 = 4'h1 == _T_88561; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_998 = 4'h2 == _T_88561; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_999 = 4'h3 == _T_88561; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1000 = 4'h4 == _T_88561; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1001 = 4'h5 == _T_88561; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1002 = 4'h6 == _T_88561; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1003 = 4'h7 == _T_88561; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1004 = 4'h8 == _T_88561; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1005 = 4'h9 == _T_88561; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1006 = 4'ha == _T_88561; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1007 = 4'hb == _T_88561; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1008 = 4'hc == _T_88561; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1009 = 4'hd == _T_88561; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1010 = 4'he == _T_88561; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1011 = 4'hf == _T_88561; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1013 = 4'h1 == _T_88561 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1014 = 4'h2 == _T_88561 ? shiftedStoreDataKnownPReg_2 : _GEN_1013; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1015 = 4'h3 == _T_88561 ? shiftedStoreDataKnownPReg_3 : _GEN_1014; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1016 = 4'h4 == _T_88561 ? shiftedStoreDataKnownPReg_4 : _GEN_1015; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1017 = 4'h5 == _T_88561 ? shiftedStoreDataKnownPReg_5 : _GEN_1016; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1018 = 4'h6 == _T_88561 ? shiftedStoreDataKnownPReg_6 : _GEN_1017; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1019 = 4'h7 == _T_88561 ? shiftedStoreDataKnownPReg_7 : _GEN_1018; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1020 = 4'h8 == _T_88561 ? shiftedStoreDataKnownPReg_8 : _GEN_1019; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1021 = 4'h9 == _T_88561 ? shiftedStoreDataKnownPReg_9 : _GEN_1020; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1022 = 4'ha == _T_88561 ? shiftedStoreDataKnownPReg_10 : _GEN_1021; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1023 = 4'hb == _T_88561 ? shiftedStoreDataKnownPReg_11 : _GEN_1022; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1024 = 4'hc == _T_88561 ? shiftedStoreDataKnownPReg_12 : _GEN_1023; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1025 = 4'hd == _T_88561 ? shiftedStoreDataKnownPReg_13 : _GEN_1024; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1026 = 4'he == _T_88561 ? shiftedStoreDataKnownPReg_14 : _GEN_1025; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1027 = 4'hf == _T_88561 ? shiftedStoreDataKnownPReg_15 : _GEN_1026; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1029 = 4'h1 == _T_88561 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1030 = 4'h2 == _T_88561 ? shiftedStoreDataQPreg_2 : _GEN_1029; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1031 = 4'h3 == _T_88561 ? shiftedStoreDataQPreg_3 : _GEN_1030; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1032 = 4'h4 == _T_88561 ? shiftedStoreDataQPreg_4 : _GEN_1031; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1033 = 4'h5 == _T_88561 ? shiftedStoreDataQPreg_5 : _GEN_1032; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1034 = 4'h6 == _T_88561 ? shiftedStoreDataQPreg_6 : _GEN_1033; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1035 = 4'h7 == _T_88561 ? shiftedStoreDataQPreg_7 : _GEN_1034; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1036 = 4'h8 == _T_88561 ? shiftedStoreDataQPreg_8 : _GEN_1035; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1037 = 4'h9 == _T_88561 ? shiftedStoreDataQPreg_9 : _GEN_1036; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1038 = 4'ha == _T_88561 ? shiftedStoreDataQPreg_10 : _GEN_1037; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1039 = 4'hb == _T_88561 ? shiftedStoreDataQPreg_11 : _GEN_1038; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1040 = 4'hc == _T_88561 ? shiftedStoreDataQPreg_12 : _GEN_1039; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1041 = 4'hd == _T_88561 ? shiftedStoreDataQPreg_13 : _GEN_1040; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1042 = 4'he == _T_88561 ? shiftedStoreDataQPreg_14 : _GEN_1041; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1043 = 4'hf == _T_88561 ? shiftedStoreDataQPreg_15 : _GEN_1042; // @[LoadQueue.scala 195:31:@35350.6]
  assign lastConflict_2_0 = _T_88578 ? _GEN_996 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_1 = _T_88578 ? _GEN_997 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_2 = _T_88578 ? _GEN_998 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_3 = _T_88578 ? _GEN_999 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_4 = _T_88578 ? _GEN_1000 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_5 = _T_88578 ? _GEN_1001 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_6 = _T_88578 ? _GEN_1002 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_7 = _T_88578 ? _GEN_1003 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_8 = _T_88578 ? _GEN_1004 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_9 = _T_88578 ? _GEN_1005 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_10 = _T_88578 ? _GEN_1006 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_11 = _T_88578 ? _GEN_1007 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_12 = _T_88578 ? _GEN_1008 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_13 = _T_88578 ? _GEN_1009 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_14 = _T_88578 ? _GEN_1010 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_15 = _T_88578 ? _GEN_1011 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign canBypass_2 = _T_88578 ? _GEN_1027 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign bypassVal_2 = _T_88578 ? _GEN_1043 : 32'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign _T_88684 = conflictPReg_3_2 ? 2'h2 : {{1'd0}, conflictPReg_3_1}; // @[LoadQueue.scala 191:60:@35404.4]
  assign _T_88685 = conflictPReg_3_3 ? 2'h3 : _T_88684; // @[LoadQueue.scala 191:60:@35405.4]
  assign _T_88686 = conflictPReg_3_4 ? 3'h4 : {{1'd0}, _T_88685}; // @[LoadQueue.scala 191:60:@35406.4]
  assign _T_88687 = conflictPReg_3_5 ? 3'h5 : _T_88686; // @[LoadQueue.scala 191:60:@35407.4]
  assign _T_88688 = conflictPReg_3_6 ? 3'h6 : _T_88687; // @[LoadQueue.scala 191:60:@35408.4]
  assign _T_88689 = conflictPReg_3_7 ? 3'h7 : _T_88688; // @[LoadQueue.scala 191:60:@35409.4]
  assign _T_88690 = conflictPReg_3_8 ? 4'h8 : {{1'd0}, _T_88689}; // @[LoadQueue.scala 191:60:@35410.4]
  assign _T_88691 = conflictPReg_3_9 ? 4'h9 : _T_88690; // @[LoadQueue.scala 191:60:@35411.4]
  assign _T_88692 = conflictPReg_3_10 ? 4'ha : _T_88691; // @[LoadQueue.scala 191:60:@35412.4]
  assign _T_88693 = conflictPReg_3_11 ? 4'hb : _T_88692; // @[LoadQueue.scala 191:60:@35413.4]
  assign _T_88694 = conflictPReg_3_12 ? 4'hc : _T_88693; // @[LoadQueue.scala 191:60:@35414.4]
  assign _T_88695 = conflictPReg_3_13 ? 4'hd : _T_88694; // @[LoadQueue.scala 191:60:@35415.4]
  assign _T_88696 = conflictPReg_3_14 ? 4'he : _T_88695; // @[LoadQueue.scala 191:60:@35416.4]
  assign _T_88697 = conflictPReg_3_15 ? 4'hf : _T_88696; // @[LoadQueue.scala 191:60:@35417.4]
  assign _T_88700 = conflictPReg_3_0 | conflictPReg_3_1; // @[LoadQueue.scala 192:43:@35419.4]
  assign _T_88701 = _T_88700 | conflictPReg_3_2; // @[LoadQueue.scala 192:43:@35420.4]
  assign _T_88702 = _T_88701 | conflictPReg_3_3; // @[LoadQueue.scala 192:43:@35421.4]
  assign _T_88703 = _T_88702 | conflictPReg_3_4; // @[LoadQueue.scala 192:43:@35422.4]
  assign _T_88704 = _T_88703 | conflictPReg_3_5; // @[LoadQueue.scala 192:43:@35423.4]
  assign _T_88705 = _T_88704 | conflictPReg_3_6; // @[LoadQueue.scala 192:43:@35424.4]
  assign _T_88706 = _T_88705 | conflictPReg_3_7; // @[LoadQueue.scala 192:43:@35425.4]
  assign _T_88707 = _T_88706 | conflictPReg_3_8; // @[LoadQueue.scala 192:43:@35426.4]
  assign _T_88708 = _T_88707 | conflictPReg_3_9; // @[LoadQueue.scala 192:43:@35427.4]
  assign _T_88709 = _T_88708 | conflictPReg_3_10; // @[LoadQueue.scala 192:43:@35428.4]
  assign _T_88710 = _T_88709 | conflictPReg_3_11; // @[LoadQueue.scala 192:43:@35429.4]
  assign _T_88711 = _T_88710 | conflictPReg_3_12; // @[LoadQueue.scala 192:43:@35430.4]
  assign _T_88712 = _T_88711 | conflictPReg_3_13; // @[LoadQueue.scala 192:43:@35431.4]
  assign _T_88713 = _T_88712 | conflictPReg_3_14; // @[LoadQueue.scala 192:43:@35432.4]
  assign _T_88714 = _T_88713 | conflictPReg_3_15; // @[LoadQueue.scala 192:43:@35433.4]
  assign _GEN_1062 = 4'h0 == _T_88697; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1063 = 4'h1 == _T_88697; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1064 = 4'h2 == _T_88697; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1065 = 4'h3 == _T_88697; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1066 = 4'h4 == _T_88697; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1067 = 4'h5 == _T_88697; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1068 = 4'h6 == _T_88697; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1069 = 4'h7 == _T_88697; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1070 = 4'h8 == _T_88697; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1071 = 4'h9 == _T_88697; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1072 = 4'ha == _T_88697; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1073 = 4'hb == _T_88697; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1074 = 4'hc == _T_88697; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1075 = 4'hd == _T_88697; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1076 = 4'he == _T_88697; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1077 = 4'hf == _T_88697; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1079 = 4'h1 == _T_88697 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1080 = 4'h2 == _T_88697 ? shiftedStoreDataKnownPReg_2 : _GEN_1079; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1081 = 4'h3 == _T_88697 ? shiftedStoreDataKnownPReg_3 : _GEN_1080; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1082 = 4'h4 == _T_88697 ? shiftedStoreDataKnownPReg_4 : _GEN_1081; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1083 = 4'h5 == _T_88697 ? shiftedStoreDataKnownPReg_5 : _GEN_1082; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1084 = 4'h6 == _T_88697 ? shiftedStoreDataKnownPReg_6 : _GEN_1083; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1085 = 4'h7 == _T_88697 ? shiftedStoreDataKnownPReg_7 : _GEN_1084; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1086 = 4'h8 == _T_88697 ? shiftedStoreDataKnownPReg_8 : _GEN_1085; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1087 = 4'h9 == _T_88697 ? shiftedStoreDataKnownPReg_9 : _GEN_1086; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1088 = 4'ha == _T_88697 ? shiftedStoreDataKnownPReg_10 : _GEN_1087; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1089 = 4'hb == _T_88697 ? shiftedStoreDataKnownPReg_11 : _GEN_1088; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1090 = 4'hc == _T_88697 ? shiftedStoreDataKnownPReg_12 : _GEN_1089; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1091 = 4'hd == _T_88697 ? shiftedStoreDataKnownPReg_13 : _GEN_1090; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1092 = 4'he == _T_88697 ? shiftedStoreDataKnownPReg_14 : _GEN_1091; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1093 = 4'hf == _T_88697 ? shiftedStoreDataKnownPReg_15 : _GEN_1092; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1095 = 4'h1 == _T_88697 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1096 = 4'h2 == _T_88697 ? shiftedStoreDataQPreg_2 : _GEN_1095; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1097 = 4'h3 == _T_88697 ? shiftedStoreDataQPreg_3 : _GEN_1096; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1098 = 4'h4 == _T_88697 ? shiftedStoreDataQPreg_4 : _GEN_1097; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1099 = 4'h5 == _T_88697 ? shiftedStoreDataQPreg_5 : _GEN_1098; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1100 = 4'h6 == _T_88697 ? shiftedStoreDataQPreg_6 : _GEN_1099; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1101 = 4'h7 == _T_88697 ? shiftedStoreDataQPreg_7 : _GEN_1100; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1102 = 4'h8 == _T_88697 ? shiftedStoreDataQPreg_8 : _GEN_1101; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1103 = 4'h9 == _T_88697 ? shiftedStoreDataQPreg_9 : _GEN_1102; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1104 = 4'ha == _T_88697 ? shiftedStoreDataQPreg_10 : _GEN_1103; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1105 = 4'hb == _T_88697 ? shiftedStoreDataQPreg_11 : _GEN_1104; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1106 = 4'hc == _T_88697 ? shiftedStoreDataQPreg_12 : _GEN_1105; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1107 = 4'hd == _T_88697 ? shiftedStoreDataQPreg_13 : _GEN_1106; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1108 = 4'he == _T_88697 ? shiftedStoreDataQPreg_14 : _GEN_1107; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1109 = 4'hf == _T_88697 ? shiftedStoreDataQPreg_15 : _GEN_1108; // @[LoadQueue.scala 195:31:@35437.6]
  assign lastConflict_3_0 = _T_88714 ? _GEN_1062 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_1 = _T_88714 ? _GEN_1063 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_2 = _T_88714 ? _GEN_1064 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_3 = _T_88714 ? _GEN_1065 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_4 = _T_88714 ? _GEN_1066 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_5 = _T_88714 ? _GEN_1067 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_6 = _T_88714 ? _GEN_1068 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_7 = _T_88714 ? _GEN_1069 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_8 = _T_88714 ? _GEN_1070 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_9 = _T_88714 ? _GEN_1071 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_10 = _T_88714 ? _GEN_1072 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_11 = _T_88714 ? _GEN_1073 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_12 = _T_88714 ? _GEN_1074 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_13 = _T_88714 ? _GEN_1075 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_14 = _T_88714 ? _GEN_1076 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_15 = _T_88714 ? _GEN_1077 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign canBypass_3 = _T_88714 ? _GEN_1093 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign bypassVal_3 = _T_88714 ? _GEN_1109 : 32'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign _T_88820 = conflictPReg_4_2 ? 2'h2 : {{1'd0}, conflictPReg_4_1}; // @[LoadQueue.scala 191:60:@35491.4]
  assign _T_88821 = conflictPReg_4_3 ? 2'h3 : _T_88820; // @[LoadQueue.scala 191:60:@35492.4]
  assign _T_88822 = conflictPReg_4_4 ? 3'h4 : {{1'd0}, _T_88821}; // @[LoadQueue.scala 191:60:@35493.4]
  assign _T_88823 = conflictPReg_4_5 ? 3'h5 : _T_88822; // @[LoadQueue.scala 191:60:@35494.4]
  assign _T_88824 = conflictPReg_4_6 ? 3'h6 : _T_88823; // @[LoadQueue.scala 191:60:@35495.4]
  assign _T_88825 = conflictPReg_4_7 ? 3'h7 : _T_88824; // @[LoadQueue.scala 191:60:@35496.4]
  assign _T_88826 = conflictPReg_4_8 ? 4'h8 : {{1'd0}, _T_88825}; // @[LoadQueue.scala 191:60:@35497.4]
  assign _T_88827 = conflictPReg_4_9 ? 4'h9 : _T_88826; // @[LoadQueue.scala 191:60:@35498.4]
  assign _T_88828 = conflictPReg_4_10 ? 4'ha : _T_88827; // @[LoadQueue.scala 191:60:@35499.4]
  assign _T_88829 = conflictPReg_4_11 ? 4'hb : _T_88828; // @[LoadQueue.scala 191:60:@35500.4]
  assign _T_88830 = conflictPReg_4_12 ? 4'hc : _T_88829; // @[LoadQueue.scala 191:60:@35501.4]
  assign _T_88831 = conflictPReg_4_13 ? 4'hd : _T_88830; // @[LoadQueue.scala 191:60:@35502.4]
  assign _T_88832 = conflictPReg_4_14 ? 4'he : _T_88831; // @[LoadQueue.scala 191:60:@35503.4]
  assign _T_88833 = conflictPReg_4_15 ? 4'hf : _T_88832; // @[LoadQueue.scala 191:60:@35504.4]
  assign _T_88836 = conflictPReg_4_0 | conflictPReg_4_1; // @[LoadQueue.scala 192:43:@35506.4]
  assign _T_88837 = _T_88836 | conflictPReg_4_2; // @[LoadQueue.scala 192:43:@35507.4]
  assign _T_88838 = _T_88837 | conflictPReg_4_3; // @[LoadQueue.scala 192:43:@35508.4]
  assign _T_88839 = _T_88838 | conflictPReg_4_4; // @[LoadQueue.scala 192:43:@35509.4]
  assign _T_88840 = _T_88839 | conflictPReg_4_5; // @[LoadQueue.scala 192:43:@35510.4]
  assign _T_88841 = _T_88840 | conflictPReg_4_6; // @[LoadQueue.scala 192:43:@35511.4]
  assign _T_88842 = _T_88841 | conflictPReg_4_7; // @[LoadQueue.scala 192:43:@35512.4]
  assign _T_88843 = _T_88842 | conflictPReg_4_8; // @[LoadQueue.scala 192:43:@35513.4]
  assign _T_88844 = _T_88843 | conflictPReg_4_9; // @[LoadQueue.scala 192:43:@35514.4]
  assign _T_88845 = _T_88844 | conflictPReg_4_10; // @[LoadQueue.scala 192:43:@35515.4]
  assign _T_88846 = _T_88845 | conflictPReg_4_11; // @[LoadQueue.scala 192:43:@35516.4]
  assign _T_88847 = _T_88846 | conflictPReg_4_12; // @[LoadQueue.scala 192:43:@35517.4]
  assign _T_88848 = _T_88847 | conflictPReg_4_13; // @[LoadQueue.scala 192:43:@35518.4]
  assign _T_88849 = _T_88848 | conflictPReg_4_14; // @[LoadQueue.scala 192:43:@35519.4]
  assign _T_88850 = _T_88849 | conflictPReg_4_15; // @[LoadQueue.scala 192:43:@35520.4]
  assign _GEN_1128 = 4'h0 == _T_88833; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1129 = 4'h1 == _T_88833; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1130 = 4'h2 == _T_88833; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1131 = 4'h3 == _T_88833; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1132 = 4'h4 == _T_88833; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1133 = 4'h5 == _T_88833; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1134 = 4'h6 == _T_88833; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1135 = 4'h7 == _T_88833; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1136 = 4'h8 == _T_88833; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1137 = 4'h9 == _T_88833; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1138 = 4'ha == _T_88833; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1139 = 4'hb == _T_88833; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1140 = 4'hc == _T_88833; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1141 = 4'hd == _T_88833; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1142 = 4'he == _T_88833; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1143 = 4'hf == _T_88833; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1145 = 4'h1 == _T_88833 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1146 = 4'h2 == _T_88833 ? shiftedStoreDataKnownPReg_2 : _GEN_1145; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1147 = 4'h3 == _T_88833 ? shiftedStoreDataKnownPReg_3 : _GEN_1146; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1148 = 4'h4 == _T_88833 ? shiftedStoreDataKnownPReg_4 : _GEN_1147; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1149 = 4'h5 == _T_88833 ? shiftedStoreDataKnownPReg_5 : _GEN_1148; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1150 = 4'h6 == _T_88833 ? shiftedStoreDataKnownPReg_6 : _GEN_1149; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1151 = 4'h7 == _T_88833 ? shiftedStoreDataKnownPReg_7 : _GEN_1150; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1152 = 4'h8 == _T_88833 ? shiftedStoreDataKnownPReg_8 : _GEN_1151; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1153 = 4'h9 == _T_88833 ? shiftedStoreDataKnownPReg_9 : _GEN_1152; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1154 = 4'ha == _T_88833 ? shiftedStoreDataKnownPReg_10 : _GEN_1153; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1155 = 4'hb == _T_88833 ? shiftedStoreDataKnownPReg_11 : _GEN_1154; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1156 = 4'hc == _T_88833 ? shiftedStoreDataKnownPReg_12 : _GEN_1155; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1157 = 4'hd == _T_88833 ? shiftedStoreDataKnownPReg_13 : _GEN_1156; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1158 = 4'he == _T_88833 ? shiftedStoreDataKnownPReg_14 : _GEN_1157; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1159 = 4'hf == _T_88833 ? shiftedStoreDataKnownPReg_15 : _GEN_1158; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1161 = 4'h1 == _T_88833 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1162 = 4'h2 == _T_88833 ? shiftedStoreDataQPreg_2 : _GEN_1161; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1163 = 4'h3 == _T_88833 ? shiftedStoreDataQPreg_3 : _GEN_1162; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1164 = 4'h4 == _T_88833 ? shiftedStoreDataQPreg_4 : _GEN_1163; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1165 = 4'h5 == _T_88833 ? shiftedStoreDataQPreg_5 : _GEN_1164; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1166 = 4'h6 == _T_88833 ? shiftedStoreDataQPreg_6 : _GEN_1165; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1167 = 4'h7 == _T_88833 ? shiftedStoreDataQPreg_7 : _GEN_1166; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1168 = 4'h8 == _T_88833 ? shiftedStoreDataQPreg_8 : _GEN_1167; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1169 = 4'h9 == _T_88833 ? shiftedStoreDataQPreg_9 : _GEN_1168; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1170 = 4'ha == _T_88833 ? shiftedStoreDataQPreg_10 : _GEN_1169; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1171 = 4'hb == _T_88833 ? shiftedStoreDataQPreg_11 : _GEN_1170; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1172 = 4'hc == _T_88833 ? shiftedStoreDataQPreg_12 : _GEN_1171; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1173 = 4'hd == _T_88833 ? shiftedStoreDataQPreg_13 : _GEN_1172; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1174 = 4'he == _T_88833 ? shiftedStoreDataQPreg_14 : _GEN_1173; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1175 = 4'hf == _T_88833 ? shiftedStoreDataQPreg_15 : _GEN_1174; // @[LoadQueue.scala 195:31:@35524.6]
  assign lastConflict_4_0 = _T_88850 ? _GEN_1128 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_1 = _T_88850 ? _GEN_1129 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_2 = _T_88850 ? _GEN_1130 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_3 = _T_88850 ? _GEN_1131 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_4 = _T_88850 ? _GEN_1132 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_5 = _T_88850 ? _GEN_1133 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_6 = _T_88850 ? _GEN_1134 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_7 = _T_88850 ? _GEN_1135 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_8 = _T_88850 ? _GEN_1136 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_9 = _T_88850 ? _GEN_1137 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_10 = _T_88850 ? _GEN_1138 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_11 = _T_88850 ? _GEN_1139 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_12 = _T_88850 ? _GEN_1140 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_13 = _T_88850 ? _GEN_1141 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_14 = _T_88850 ? _GEN_1142 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_15 = _T_88850 ? _GEN_1143 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign canBypass_4 = _T_88850 ? _GEN_1159 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign bypassVal_4 = _T_88850 ? _GEN_1175 : 32'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign _T_88956 = conflictPReg_5_2 ? 2'h2 : {{1'd0}, conflictPReg_5_1}; // @[LoadQueue.scala 191:60:@35578.4]
  assign _T_88957 = conflictPReg_5_3 ? 2'h3 : _T_88956; // @[LoadQueue.scala 191:60:@35579.4]
  assign _T_88958 = conflictPReg_5_4 ? 3'h4 : {{1'd0}, _T_88957}; // @[LoadQueue.scala 191:60:@35580.4]
  assign _T_88959 = conflictPReg_5_5 ? 3'h5 : _T_88958; // @[LoadQueue.scala 191:60:@35581.4]
  assign _T_88960 = conflictPReg_5_6 ? 3'h6 : _T_88959; // @[LoadQueue.scala 191:60:@35582.4]
  assign _T_88961 = conflictPReg_5_7 ? 3'h7 : _T_88960; // @[LoadQueue.scala 191:60:@35583.4]
  assign _T_88962 = conflictPReg_5_8 ? 4'h8 : {{1'd0}, _T_88961}; // @[LoadQueue.scala 191:60:@35584.4]
  assign _T_88963 = conflictPReg_5_9 ? 4'h9 : _T_88962; // @[LoadQueue.scala 191:60:@35585.4]
  assign _T_88964 = conflictPReg_5_10 ? 4'ha : _T_88963; // @[LoadQueue.scala 191:60:@35586.4]
  assign _T_88965 = conflictPReg_5_11 ? 4'hb : _T_88964; // @[LoadQueue.scala 191:60:@35587.4]
  assign _T_88966 = conflictPReg_5_12 ? 4'hc : _T_88965; // @[LoadQueue.scala 191:60:@35588.4]
  assign _T_88967 = conflictPReg_5_13 ? 4'hd : _T_88966; // @[LoadQueue.scala 191:60:@35589.4]
  assign _T_88968 = conflictPReg_5_14 ? 4'he : _T_88967; // @[LoadQueue.scala 191:60:@35590.4]
  assign _T_88969 = conflictPReg_5_15 ? 4'hf : _T_88968; // @[LoadQueue.scala 191:60:@35591.4]
  assign _T_88972 = conflictPReg_5_0 | conflictPReg_5_1; // @[LoadQueue.scala 192:43:@35593.4]
  assign _T_88973 = _T_88972 | conflictPReg_5_2; // @[LoadQueue.scala 192:43:@35594.4]
  assign _T_88974 = _T_88973 | conflictPReg_5_3; // @[LoadQueue.scala 192:43:@35595.4]
  assign _T_88975 = _T_88974 | conflictPReg_5_4; // @[LoadQueue.scala 192:43:@35596.4]
  assign _T_88976 = _T_88975 | conflictPReg_5_5; // @[LoadQueue.scala 192:43:@35597.4]
  assign _T_88977 = _T_88976 | conflictPReg_5_6; // @[LoadQueue.scala 192:43:@35598.4]
  assign _T_88978 = _T_88977 | conflictPReg_5_7; // @[LoadQueue.scala 192:43:@35599.4]
  assign _T_88979 = _T_88978 | conflictPReg_5_8; // @[LoadQueue.scala 192:43:@35600.4]
  assign _T_88980 = _T_88979 | conflictPReg_5_9; // @[LoadQueue.scala 192:43:@35601.4]
  assign _T_88981 = _T_88980 | conflictPReg_5_10; // @[LoadQueue.scala 192:43:@35602.4]
  assign _T_88982 = _T_88981 | conflictPReg_5_11; // @[LoadQueue.scala 192:43:@35603.4]
  assign _T_88983 = _T_88982 | conflictPReg_5_12; // @[LoadQueue.scala 192:43:@35604.4]
  assign _T_88984 = _T_88983 | conflictPReg_5_13; // @[LoadQueue.scala 192:43:@35605.4]
  assign _T_88985 = _T_88984 | conflictPReg_5_14; // @[LoadQueue.scala 192:43:@35606.4]
  assign _T_88986 = _T_88985 | conflictPReg_5_15; // @[LoadQueue.scala 192:43:@35607.4]
  assign _GEN_1194 = 4'h0 == _T_88969; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1195 = 4'h1 == _T_88969; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1196 = 4'h2 == _T_88969; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1197 = 4'h3 == _T_88969; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1198 = 4'h4 == _T_88969; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1199 = 4'h5 == _T_88969; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1200 = 4'h6 == _T_88969; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1201 = 4'h7 == _T_88969; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1202 = 4'h8 == _T_88969; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1203 = 4'h9 == _T_88969; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1204 = 4'ha == _T_88969; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1205 = 4'hb == _T_88969; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1206 = 4'hc == _T_88969; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1207 = 4'hd == _T_88969; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1208 = 4'he == _T_88969; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1209 = 4'hf == _T_88969; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1211 = 4'h1 == _T_88969 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1212 = 4'h2 == _T_88969 ? shiftedStoreDataKnownPReg_2 : _GEN_1211; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1213 = 4'h3 == _T_88969 ? shiftedStoreDataKnownPReg_3 : _GEN_1212; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1214 = 4'h4 == _T_88969 ? shiftedStoreDataKnownPReg_4 : _GEN_1213; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1215 = 4'h5 == _T_88969 ? shiftedStoreDataKnownPReg_5 : _GEN_1214; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1216 = 4'h6 == _T_88969 ? shiftedStoreDataKnownPReg_6 : _GEN_1215; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1217 = 4'h7 == _T_88969 ? shiftedStoreDataKnownPReg_7 : _GEN_1216; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1218 = 4'h8 == _T_88969 ? shiftedStoreDataKnownPReg_8 : _GEN_1217; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1219 = 4'h9 == _T_88969 ? shiftedStoreDataKnownPReg_9 : _GEN_1218; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1220 = 4'ha == _T_88969 ? shiftedStoreDataKnownPReg_10 : _GEN_1219; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1221 = 4'hb == _T_88969 ? shiftedStoreDataKnownPReg_11 : _GEN_1220; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1222 = 4'hc == _T_88969 ? shiftedStoreDataKnownPReg_12 : _GEN_1221; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1223 = 4'hd == _T_88969 ? shiftedStoreDataKnownPReg_13 : _GEN_1222; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1224 = 4'he == _T_88969 ? shiftedStoreDataKnownPReg_14 : _GEN_1223; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1225 = 4'hf == _T_88969 ? shiftedStoreDataKnownPReg_15 : _GEN_1224; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1227 = 4'h1 == _T_88969 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1228 = 4'h2 == _T_88969 ? shiftedStoreDataQPreg_2 : _GEN_1227; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1229 = 4'h3 == _T_88969 ? shiftedStoreDataQPreg_3 : _GEN_1228; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1230 = 4'h4 == _T_88969 ? shiftedStoreDataQPreg_4 : _GEN_1229; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1231 = 4'h5 == _T_88969 ? shiftedStoreDataQPreg_5 : _GEN_1230; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1232 = 4'h6 == _T_88969 ? shiftedStoreDataQPreg_6 : _GEN_1231; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1233 = 4'h7 == _T_88969 ? shiftedStoreDataQPreg_7 : _GEN_1232; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1234 = 4'h8 == _T_88969 ? shiftedStoreDataQPreg_8 : _GEN_1233; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1235 = 4'h9 == _T_88969 ? shiftedStoreDataQPreg_9 : _GEN_1234; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1236 = 4'ha == _T_88969 ? shiftedStoreDataQPreg_10 : _GEN_1235; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1237 = 4'hb == _T_88969 ? shiftedStoreDataQPreg_11 : _GEN_1236; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1238 = 4'hc == _T_88969 ? shiftedStoreDataQPreg_12 : _GEN_1237; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1239 = 4'hd == _T_88969 ? shiftedStoreDataQPreg_13 : _GEN_1238; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1240 = 4'he == _T_88969 ? shiftedStoreDataQPreg_14 : _GEN_1239; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1241 = 4'hf == _T_88969 ? shiftedStoreDataQPreg_15 : _GEN_1240; // @[LoadQueue.scala 195:31:@35611.6]
  assign lastConflict_5_0 = _T_88986 ? _GEN_1194 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_1 = _T_88986 ? _GEN_1195 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_2 = _T_88986 ? _GEN_1196 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_3 = _T_88986 ? _GEN_1197 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_4 = _T_88986 ? _GEN_1198 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_5 = _T_88986 ? _GEN_1199 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_6 = _T_88986 ? _GEN_1200 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_7 = _T_88986 ? _GEN_1201 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_8 = _T_88986 ? _GEN_1202 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_9 = _T_88986 ? _GEN_1203 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_10 = _T_88986 ? _GEN_1204 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_11 = _T_88986 ? _GEN_1205 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_12 = _T_88986 ? _GEN_1206 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_13 = _T_88986 ? _GEN_1207 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_14 = _T_88986 ? _GEN_1208 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_15 = _T_88986 ? _GEN_1209 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign canBypass_5 = _T_88986 ? _GEN_1225 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign bypassVal_5 = _T_88986 ? _GEN_1241 : 32'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign _T_89092 = conflictPReg_6_2 ? 2'h2 : {{1'd0}, conflictPReg_6_1}; // @[LoadQueue.scala 191:60:@35665.4]
  assign _T_89093 = conflictPReg_6_3 ? 2'h3 : _T_89092; // @[LoadQueue.scala 191:60:@35666.4]
  assign _T_89094 = conflictPReg_6_4 ? 3'h4 : {{1'd0}, _T_89093}; // @[LoadQueue.scala 191:60:@35667.4]
  assign _T_89095 = conflictPReg_6_5 ? 3'h5 : _T_89094; // @[LoadQueue.scala 191:60:@35668.4]
  assign _T_89096 = conflictPReg_6_6 ? 3'h6 : _T_89095; // @[LoadQueue.scala 191:60:@35669.4]
  assign _T_89097 = conflictPReg_6_7 ? 3'h7 : _T_89096; // @[LoadQueue.scala 191:60:@35670.4]
  assign _T_89098 = conflictPReg_6_8 ? 4'h8 : {{1'd0}, _T_89097}; // @[LoadQueue.scala 191:60:@35671.4]
  assign _T_89099 = conflictPReg_6_9 ? 4'h9 : _T_89098; // @[LoadQueue.scala 191:60:@35672.4]
  assign _T_89100 = conflictPReg_6_10 ? 4'ha : _T_89099; // @[LoadQueue.scala 191:60:@35673.4]
  assign _T_89101 = conflictPReg_6_11 ? 4'hb : _T_89100; // @[LoadQueue.scala 191:60:@35674.4]
  assign _T_89102 = conflictPReg_6_12 ? 4'hc : _T_89101; // @[LoadQueue.scala 191:60:@35675.4]
  assign _T_89103 = conflictPReg_6_13 ? 4'hd : _T_89102; // @[LoadQueue.scala 191:60:@35676.4]
  assign _T_89104 = conflictPReg_6_14 ? 4'he : _T_89103; // @[LoadQueue.scala 191:60:@35677.4]
  assign _T_89105 = conflictPReg_6_15 ? 4'hf : _T_89104; // @[LoadQueue.scala 191:60:@35678.4]
  assign _T_89108 = conflictPReg_6_0 | conflictPReg_6_1; // @[LoadQueue.scala 192:43:@35680.4]
  assign _T_89109 = _T_89108 | conflictPReg_6_2; // @[LoadQueue.scala 192:43:@35681.4]
  assign _T_89110 = _T_89109 | conflictPReg_6_3; // @[LoadQueue.scala 192:43:@35682.4]
  assign _T_89111 = _T_89110 | conflictPReg_6_4; // @[LoadQueue.scala 192:43:@35683.4]
  assign _T_89112 = _T_89111 | conflictPReg_6_5; // @[LoadQueue.scala 192:43:@35684.4]
  assign _T_89113 = _T_89112 | conflictPReg_6_6; // @[LoadQueue.scala 192:43:@35685.4]
  assign _T_89114 = _T_89113 | conflictPReg_6_7; // @[LoadQueue.scala 192:43:@35686.4]
  assign _T_89115 = _T_89114 | conflictPReg_6_8; // @[LoadQueue.scala 192:43:@35687.4]
  assign _T_89116 = _T_89115 | conflictPReg_6_9; // @[LoadQueue.scala 192:43:@35688.4]
  assign _T_89117 = _T_89116 | conflictPReg_6_10; // @[LoadQueue.scala 192:43:@35689.4]
  assign _T_89118 = _T_89117 | conflictPReg_6_11; // @[LoadQueue.scala 192:43:@35690.4]
  assign _T_89119 = _T_89118 | conflictPReg_6_12; // @[LoadQueue.scala 192:43:@35691.4]
  assign _T_89120 = _T_89119 | conflictPReg_6_13; // @[LoadQueue.scala 192:43:@35692.4]
  assign _T_89121 = _T_89120 | conflictPReg_6_14; // @[LoadQueue.scala 192:43:@35693.4]
  assign _T_89122 = _T_89121 | conflictPReg_6_15; // @[LoadQueue.scala 192:43:@35694.4]
  assign _GEN_1260 = 4'h0 == _T_89105; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1261 = 4'h1 == _T_89105; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1262 = 4'h2 == _T_89105; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1263 = 4'h3 == _T_89105; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1264 = 4'h4 == _T_89105; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1265 = 4'h5 == _T_89105; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1266 = 4'h6 == _T_89105; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1267 = 4'h7 == _T_89105; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1268 = 4'h8 == _T_89105; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1269 = 4'h9 == _T_89105; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1270 = 4'ha == _T_89105; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1271 = 4'hb == _T_89105; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1272 = 4'hc == _T_89105; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1273 = 4'hd == _T_89105; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1274 = 4'he == _T_89105; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1275 = 4'hf == _T_89105; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1277 = 4'h1 == _T_89105 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1278 = 4'h2 == _T_89105 ? shiftedStoreDataKnownPReg_2 : _GEN_1277; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1279 = 4'h3 == _T_89105 ? shiftedStoreDataKnownPReg_3 : _GEN_1278; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1280 = 4'h4 == _T_89105 ? shiftedStoreDataKnownPReg_4 : _GEN_1279; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1281 = 4'h5 == _T_89105 ? shiftedStoreDataKnownPReg_5 : _GEN_1280; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1282 = 4'h6 == _T_89105 ? shiftedStoreDataKnownPReg_6 : _GEN_1281; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1283 = 4'h7 == _T_89105 ? shiftedStoreDataKnownPReg_7 : _GEN_1282; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1284 = 4'h8 == _T_89105 ? shiftedStoreDataKnownPReg_8 : _GEN_1283; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1285 = 4'h9 == _T_89105 ? shiftedStoreDataKnownPReg_9 : _GEN_1284; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1286 = 4'ha == _T_89105 ? shiftedStoreDataKnownPReg_10 : _GEN_1285; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1287 = 4'hb == _T_89105 ? shiftedStoreDataKnownPReg_11 : _GEN_1286; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1288 = 4'hc == _T_89105 ? shiftedStoreDataKnownPReg_12 : _GEN_1287; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1289 = 4'hd == _T_89105 ? shiftedStoreDataKnownPReg_13 : _GEN_1288; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1290 = 4'he == _T_89105 ? shiftedStoreDataKnownPReg_14 : _GEN_1289; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1291 = 4'hf == _T_89105 ? shiftedStoreDataKnownPReg_15 : _GEN_1290; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1293 = 4'h1 == _T_89105 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1294 = 4'h2 == _T_89105 ? shiftedStoreDataQPreg_2 : _GEN_1293; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1295 = 4'h3 == _T_89105 ? shiftedStoreDataQPreg_3 : _GEN_1294; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1296 = 4'h4 == _T_89105 ? shiftedStoreDataQPreg_4 : _GEN_1295; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1297 = 4'h5 == _T_89105 ? shiftedStoreDataQPreg_5 : _GEN_1296; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1298 = 4'h6 == _T_89105 ? shiftedStoreDataQPreg_6 : _GEN_1297; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1299 = 4'h7 == _T_89105 ? shiftedStoreDataQPreg_7 : _GEN_1298; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1300 = 4'h8 == _T_89105 ? shiftedStoreDataQPreg_8 : _GEN_1299; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1301 = 4'h9 == _T_89105 ? shiftedStoreDataQPreg_9 : _GEN_1300; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1302 = 4'ha == _T_89105 ? shiftedStoreDataQPreg_10 : _GEN_1301; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1303 = 4'hb == _T_89105 ? shiftedStoreDataQPreg_11 : _GEN_1302; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1304 = 4'hc == _T_89105 ? shiftedStoreDataQPreg_12 : _GEN_1303; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1305 = 4'hd == _T_89105 ? shiftedStoreDataQPreg_13 : _GEN_1304; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1306 = 4'he == _T_89105 ? shiftedStoreDataQPreg_14 : _GEN_1305; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1307 = 4'hf == _T_89105 ? shiftedStoreDataQPreg_15 : _GEN_1306; // @[LoadQueue.scala 195:31:@35698.6]
  assign lastConflict_6_0 = _T_89122 ? _GEN_1260 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_1 = _T_89122 ? _GEN_1261 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_2 = _T_89122 ? _GEN_1262 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_3 = _T_89122 ? _GEN_1263 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_4 = _T_89122 ? _GEN_1264 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_5 = _T_89122 ? _GEN_1265 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_6 = _T_89122 ? _GEN_1266 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_7 = _T_89122 ? _GEN_1267 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_8 = _T_89122 ? _GEN_1268 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_9 = _T_89122 ? _GEN_1269 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_10 = _T_89122 ? _GEN_1270 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_11 = _T_89122 ? _GEN_1271 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_12 = _T_89122 ? _GEN_1272 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_13 = _T_89122 ? _GEN_1273 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_14 = _T_89122 ? _GEN_1274 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_15 = _T_89122 ? _GEN_1275 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign canBypass_6 = _T_89122 ? _GEN_1291 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign bypassVal_6 = _T_89122 ? _GEN_1307 : 32'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign _T_89228 = conflictPReg_7_2 ? 2'h2 : {{1'd0}, conflictPReg_7_1}; // @[LoadQueue.scala 191:60:@35752.4]
  assign _T_89229 = conflictPReg_7_3 ? 2'h3 : _T_89228; // @[LoadQueue.scala 191:60:@35753.4]
  assign _T_89230 = conflictPReg_7_4 ? 3'h4 : {{1'd0}, _T_89229}; // @[LoadQueue.scala 191:60:@35754.4]
  assign _T_89231 = conflictPReg_7_5 ? 3'h5 : _T_89230; // @[LoadQueue.scala 191:60:@35755.4]
  assign _T_89232 = conflictPReg_7_6 ? 3'h6 : _T_89231; // @[LoadQueue.scala 191:60:@35756.4]
  assign _T_89233 = conflictPReg_7_7 ? 3'h7 : _T_89232; // @[LoadQueue.scala 191:60:@35757.4]
  assign _T_89234 = conflictPReg_7_8 ? 4'h8 : {{1'd0}, _T_89233}; // @[LoadQueue.scala 191:60:@35758.4]
  assign _T_89235 = conflictPReg_7_9 ? 4'h9 : _T_89234; // @[LoadQueue.scala 191:60:@35759.4]
  assign _T_89236 = conflictPReg_7_10 ? 4'ha : _T_89235; // @[LoadQueue.scala 191:60:@35760.4]
  assign _T_89237 = conflictPReg_7_11 ? 4'hb : _T_89236; // @[LoadQueue.scala 191:60:@35761.4]
  assign _T_89238 = conflictPReg_7_12 ? 4'hc : _T_89237; // @[LoadQueue.scala 191:60:@35762.4]
  assign _T_89239 = conflictPReg_7_13 ? 4'hd : _T_89238; // @[LoadQueue.scala 191:60:@35763.4]
  assign _T_89240 = conflictPReg_7_14 ? 4'he : _T_89239; // @[LoadQueue.scala 191:60:@35764.4]
  assign _T_89241 = conflictPReg_7_15 ? 4'hf : _T_89240; // @[LoadQueue.scala 191:60:@35765.4]
  assign _T_89244 = conflictPReg_7_0 | conflictPReg_7_1; // @[LoadQueue.scala 192:43:@35767.4]
  assign _T_89245 = _T_89244 | conflictPReg_7_2; // @[LoadQueue.scala 192:43:@35768.4]
  assign _T_89246 = _T_89245 | conflictPReg_7_3; // @[LoadQueue.scala 192:43:@35769.4]
  assign _T_89247 = _T_89246 | conflictPReg_7_4; // @[LoadQueue.scala 192:43:@35770.4]
  assign _T_89248 = _T_89247 | conflictPReg_7_5; // @[LoadQueue.scala 192:43:@35771.4]
  assign _T_89249 = _T_89248 | conflictPReg_7_6; // @[LoadQueue.scala 192:43:@35772.4]
  assign _T_89250 = _T_89249 | conflictPReg_7_7; // @[LoadQueue.scala 192:43:@35773.4]
  assign _T_89251 = _T_89250 | conflictPReg_7_8; // @[LoadQueue.scala 192:43:@35774.4]
  assign _T_89252 = _T_89251 | conflictPReg_7_9; // @[LoadQueue.scala 192:43:@35775.4]
  assign _T_89253 = _T_89252 | conflictPReg_7_10; // @[LoadQueue.scala 192:43:@35776.4]
  assign _T_89254 = _T_89253 | conflictPReg_7_11; // @[LoadQueue.scala 192:43:@35777.4]
  assign _T_89255 = _T_89254 | conflictPReg_7_12; // @[LoadQueue.scala 192:43:@35778.4]
  assign _T_89256 = _T_89255 | conflictPReg_7_13; // @[LoadQueue.scala 192:43:@35779.4]
  assign _T_89257 = _T_89256 | conflictPReg_7_14; // @[LoadQueue.scala 192:43:@35780.4]
  assign _T_89258 = _T_89257 | conflictPReg_7_15; // @[LoadQueue.scala 192:43:@35781.4]
  assign _GEN_1326 = 4'h0 == _T_89241; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1327 = 4'h1 == _T_89241; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1328 = 4'h2 == _T_89241; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1329 = 4'h3 == _T_89241; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1330 = 4'h4 == _T_89241; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1331 = 4'h5 == _T_89241; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1332 = 4'h6 == _T_89241; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1333 = 4'h7 == _T_89241; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1334 = 4'h8 == _T_89241; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1335 = 4'h9 == _T_89241; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1336 = 4'ha == _T_89241; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1337 = 4'hb == _T_89241; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1338 = 4'hc == _T_89241; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1339 = 4'hd == _T_89241; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1340 = 4'he == _T_89241; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1341 = 4'hf == _T_89241; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1343 = 4'h1 == _T_89241 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1344 = 4'h2 == _T_89241 ? shiftedStoreDataKnownPReg_2 : _GEN_1343; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1345 = 4'h3 == _T_89241 ? shiftedStoreDataKnownPReg_3 : _GEN_1344; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1346 = 4'h4 == _T_89241 ? shiftedStoreDataKnownPReg_4 : _GEN_1345; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1347 = 4'h5 == _T_89241 ? shiftedStoreDataKnownPReg_5 : _GEN_1346; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1348 = 4'h6 == _T_89241 ? shiftedStoreDataKnownPReg_6 : _GEN_1347; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1349 = 4'h7 == _T_89241 ? shiftedStoreDataKnownPReg_7 : _GEN_1348; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1350 = 4'h8 == _T_89241 ? shiftedStoreDataKnownPReg_8 : _GEN_1349; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1351 = 4'h9 == _T_89241 ? shiftedStoreDataKnownPReg_9 : _GEN_1350; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1352 = 4'ha == _T_89241 ? shiftedStoreDataKnownPReg_10 : _GEN_1351; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1353 = 4'hb == _T_89241 ? shiftedStoreDataKnownPReg_11 : _GEN_1352; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1354 = 4'hc == _T_89241 ? shiftedStoreDataKnownPReg_12 : _GEN_1353; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1355 = 4'hd == _T_89241 ? shiftedStoreDataKnownPReg_13 : _GEN_1354; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1356 = 4'he == _T_89241 ? shiftedStoreDataKnownPReg_14 : _GEN_1355; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1357 = 4'hf == _T_89241 ? shiftedStoreDataKnownPReg_15 : _GEN_1356; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1359 = 4'h1 == _T_89241 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1360 = 4'h2 == _T_89241 ? shiftedStoreDataQPreg_2 : _GEN_1359; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1361 = 4'h3 == _T_89241 ? shiftedStoreDataQPreg_3 : _GEN_1360; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1362 = 4'h4 == _T_89241 ? shiftedStoreDataQPreg_4 : _GEN_1361; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1363 = 4'h5 == _T_89241 ? shiftedStoreDataQPreg_5 : _GEN_1362; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1364 = 4'h6 == _T_89241 ? shiftedStoreDataQPreg_6 : _GEN_1363; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1365 = 4'h7 == _T_89241 ? shiftedStoreDataQPreg_7 : _GEN_1364; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1366 = 4'h8 == _T_89241 ? shiftedStoreDataQPreg_8 : _GEN_1365; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1367 = 4'h9 == _T_89241 ? shiftedStoreDataQPreg_9 : _GEN_1366; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1368 = 4'ha == _T_89241 ? shiftedStoreDataQPreg_10 : _GEN_1367; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1369 = 4'hb == _T_89241 ? shiftedStoreDataQPreg_11 : _GEN_1368; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1370 = 4'hc == _T_89241 ? shiftedStoreDataQPreg_12 : _GEN_1369; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1371 = 4'hd == _T_89241 ? shiftedStoreDataQPreg_13 : _GEN_1370; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1372 = 4'he == _T_89241 ? shiftedStoreDataQPreg_14 : _GEN_1371; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1373 = 4'hf == _T_89241 ? shiftedStoreDataQPreg_15 : _GEN_1372; // @[LoadQueue.scala 195:31:@35785.6]
  assign lastConflict_7_0 = _T_89258 ? _GEN_1326 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_1 = _T_89258 ? _GEN_1327 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_2 = _T_89258 ? _GEN_1328 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_3 = _T_89258 ? _GEN_1329 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_4 = _T_89258 ? _GEN_1330 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_5 = _T_89258 ? _GEN_1331 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_6 = _T_89258 ? _GEN_1332 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_7 = _T_89258 ? _GEN_1333 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_8 = _T_89258 ? _GEN_1334 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_9 = _T_89258 ? _GEN_1335 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_10 = _T_89258 ? _GEN_1336 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_11 = _T_89258 ? _GEN_1337 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_12 = _T_89258 ? _GEN_1338 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_13 = _T_89258 ? _GEN_1339 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_14 = _T_89258 ? _GEN_1340 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_15 = _T_89258 ? _GEN_1341 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign canBypass_7 = _T_89258 ? _GEN_1357 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign bypassVal_7 = _T_89258 ? _GEN_1373 : 32'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign _T_89364 = conflictPReg_8_2 ? 2'h2 : {{1'd0}, conflictPReg_8_1}; // @[LoadQueue.scala 191:60:@35839.4]
  assign _T_89365 = conflictPReg_8_3 ? 2'h3 : _T_89364; // @[LoadQueue.scala 191:60:@35840.4]
  assign _T_89366 = conflictPReg_8_4 ? 3'h4 : {{1'd0}, _T_89365}; // @[LoadQueue.scala 191:60:@35841.4]
  assign _T_89367 = conflictPReg_8_5 ? 3'h5 : _T_89366; // @[LoadQueue.scala 191:60:@35842.4]
  assign _T_89368 = conflictPReg_8_6 ? 3'h6 : _T_89367; // @[LoadQueue.scala 191:60:@35843.4]
  assign _T_89369 = conflictPReg_8_7 ? 3'h7 : _T_89368; // @[LoadQueue.scala 191:60:@35844.4]
  assign _T_89370 = conflictPReg_8_8 ? 4'h8 : {{1'd0}, _T_89369}; // @[LoadQueue.scala 191:60:@35845.4]
  assign _T_89371 = conflictPReg_8_9 ? 4'h9 : _T_89370; // @[LoadQueue.scala 191:60:@35846.4]
  assign _T_89372 = conflictPReg_8_10 ? 4'ha : _T_89371; // @[LoadQueue.scala 191:60:@35847.4]
  assign _T_89373 = conflictPReg_8_11 ? 4'hb : _T_89372; // @[LoadQueue.scala 191:60:@35848.4]
  assign _T_89374 = conflictPReg_8_12 ? 4'hc : _T_89373; // @[LoadQueue.scala 191:60:@35849.4]
  assign _T_89375 = conflictPReg_8_13 ? 4'hd : _T_89374; // @[LoadQueue.scala 191:60:@35850.4]
  assign _T_89376 = conflictPReg_8_14 ? 4'he : _T_89375; // @[LoadQueue.scala 191:60:@35851.4]
  assign _T_89377 = conflictPReg_8_15 ? 4'hf : _T_89376; // @[LoadQueue.scala 191:60:@35852.4]
  assign _T_89380 = conflictPReg_8_0 | conflictPReg_8_1; // @[LoadQueue.scala 192:43:@35854.4]
  assign _T_89381 = _T_89380 | conflictPReg_8_2; // @[LoadQueue.scala 192:43:@35855.4]
  assign _T_89382 = _T_89381 | conflictPReg_8_3; // @[LoadQueue.scala 192:43:@35856.4]
  assign _T_89383 = _T_89382 | conflictPReg_8_4; // @[LoadQueue.scala 192:43:@35857.4]
  assign _T_89384 = _T_89383 | conflictPReg_8_5; // @[LoadQueue.scala 192:43:@35858.4]
  assign _T_89385 = _T_89384 | conflictPReg_8_6; // @[LoadQueue.scala 192:43:@35859.4]
  assign _T_89386 = _T_89385 | conflictPReg_8_7; // @[LoadQueue.scala 192:43:@35860.4]
  assign _T_89387 = _T_89386 | conflictPReg_8_8; // @[LoadQueue.scala 192:43:@35861.4]
  assign _T_89388 = _T_89387 | conflictPReg_8_9; // @[LoadQueue.scala 192:43:@35862.4]
  assign _T_89389 = _T_89388 | conflictPReg_8_10; // @[LoadQueue.scala 192:43:@35863.4]
  assign _T_89390 = _T_89389 | conflictPReg_8_11; // @[LoadQueue.scala 192:43:@35864.4]
  assign _T_89391 = _T_89390 | conflictPReg_8_12; // @[LoadQueue.scala 192:43:@35865.4]
  assign _T_89392 = _T_89391 | conflictPReg_8_13; // @[LoadQueue.scala 192:43:@35866.4]
  assign _T_89393 = _T_89392 | conflictPReg_8_14; // @[LoadQueue.scala 192:43:@35867.4]
  assign _T_89394 = _T_89393 | conflictPReg_8_15; // @[LoadQueue.scala 192:43:@35868.4]
  assign _GEN_1392 = 4'h0 == _T_89377; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1393 = 4'h1 == _T_89377; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1394 = 4'h2 == _T_89377; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1395 = 4'h3 == _T_89377; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1396 = 4'h4 == _T_89377; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1397 = 4'h5 == _T_89377; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1398 = 4'h6 == _T_89377; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1399 = 4'h7 == _T_89377; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1400 = 4'h8 == _T_89377; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1401 = 4'h9 == _T_89377; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1402 = 4'ha == _T_89377; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1403 = 4'hb == _T_89377; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1404 = 4'hc == _T_89377; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1405 = 4'hd == _T_89377; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1406 = 4'he == _T_89377; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1407 = 4'hf == _T_89377; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1409 = 4'h1 == _T_89377 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1410 = 4'h2 == _T_89377 ? shiftedStoreDataKnownPReg_2 : _GEN_1409; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1411 = 4'h3 == _T_89377 ? shiftedStoreDataKnownPReg_3 : _GEN_1410; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1412 = 4'h4 == _T_89377 ? shiftedStoreDataKnownPReg_4 : _GEN_1411; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1413 = 4'h5 == _T_89377 ? shiftedStoreDataKnownPReg_5 : _GEN_1412; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1414 = 4'h6 == _T_89377 ? shiftedStoreDataKnownPReg_6 : _GEN_1413; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1415 = 4'h7 == _T_89377 ? shiftedStoreDataKnownPReg_7 : _GEN_1414; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1416 = 4'h8 == _T_89377 ? shiftedStoreDataKnownPReg_8 : _GEN_1415; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1417 = 4'h9 == _T_89377 ? shiftedStoreDataKnownPReg_9 : _GEN_1416; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1418 = 4'ha == _T_89377 ? shiftedStoreDataKnownPReg_10 : _GEN_1417; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1419 = 4'hb == _T_89377 ? shiftedStoreDataKnownPReg_11 : _GEN_1418; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1420 = 4'hc == _T_89377 ? shiftedStoreDataKnownPReg_12 : _GEN_1419; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1421 = 4'hd == _T_89377 ? shiftedStoreDataKnownPReg_13 : _GEN_1420; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1422 = 4'he == _T_89377 ? shiftedStoreDataKnownPReg_14 : _GEN_1421; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1423 = 4'hf == _T_89377 ? shiftedStoreDataKnownPReg_15 : _GEN_1422; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1425 = 4'h1 == _T_89377 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1426 = 4'h2 == _T_89377 ? shiftedStoreDataQPreg_2 : _GEN_1425; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1427 = 4'h3 == _T_89377 ? shiftedStoreDataQPreg_3 : _GEN_1426; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1428 = 4'h4 == _T_89377 ? shiftedStoreDataQPreg_4 : _GEN_1427; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1429 = 4'h5 == _T_89377 ? shiftedStoreDataQPreg_5 : _GEN_1428; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1430 = 4'h6 == _T_89377 ? shiftedStoreDataQPreg_6 : _GEN_1429; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1431 = 4'h7 == _T_89377 ? shiftedStoreDataQPreg_7 : _GEN_1430; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1432 = 4'h8 == _T_89377 ? shiftedStoreDataQPreg_8 : _GEN_1431; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1433 = 4'h9 == _T_89377 ? shiftedStoreDataQPreg_9 : _GEN_1432; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1434 = 4'ha == _T_89377 ? shiftedStoreDataQPreg_10 : _GEN_1433; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1435 = 4'hb == _T_89377 ? shiftedStoreDataQPreg_11 : _GEN_1434; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1436 = 4'hc == _T_89377 ? shiftedStoreDataQPreg_12 : _GEN_1435; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1437 = 4'hd == _T_89377 ? shiftedStoreDataQPreg_13 : _GEN_1436; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1438 = 4'he == _T_89377 ? shiftedStoreDataQPreg_14 : _GEN_1437; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1439 = 4'hf == _T_89377 ? shiftedStoreDataQPreg_15 : _GEN_1438; // @[LoadQueue.scala 195:31:@35872.6]
  assign lastConflict_8_0 = _T_89394 ? _GEN_1392 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_1 = _T_89394 ? _GEN_1393 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_2 = _T_89394 ? _GEN_1394 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_3 = _T_89394 ? _GEN_1395 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_4 = _T_89394 ? _GEN_1396 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_5 = _T_89394 ? _GEN_1397 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_6 = _T_89394 ? _GEN_1398 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_7 = _T_89394 ? _GEN_1399 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_8 = _T_89394 ? _GEN_1400 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_9 = _T_89394 ? _GEN_1401 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_10 = _T_89394 ? _GEN_1402 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_11 = _T_89394 ? _GEN_1403 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_12 = _T_89394 ? _GEN_1404 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_13 = _T_89394 ? _GEN_1405 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_14 = _T_89394 ? _GEN_1406 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_15 = _T_89394 ? _GEN_1407 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign canBypass_8 = _T_89394 ? _GEN_1423 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign bypassVal_8 = _T_89394 ? _GEN_1439 : 32'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign _T_89500 = conflictPReg_9_2 ? 2'h2 : {{1'd0}, conflictPReg_9_1}; // @[LoadQueue.scala 191:60:@35926.4]
  assign _T_89501 = conflictPReg_9_3 ? 2'h3 : _T_89500; // @[LoadQueue.scala 191:60:@35927.4]
  assign _T_89502 = conflictPReg_9_4 ? 3'h4 : {{1'd0}, _T_89501}; // @[LoadQueue.scala 191:60:@35928.4]
  assign _T_89503 = conflictPReg_9_5 ? 3'h5 : _T_89502; // @[LoadQueue.scala 191:60:@35929.4]
  assign _T_89504 = conflictPReg_9_6 ? 3'h6 : _T_89503; // @[LoadQueue.scala 191:60:@35930.4]
  assign _T_89505 = conflictPReg_9_7 ? 3'h7 : _T_89504; // @[LoadQueue.scala 191:60:@35931.4]
  assign _T_89506 = conflictPReg_9_8 ? 4'h8 : {{1'd0}, _T_89505}; // @[LoadQueue.scala 191:60:@35932.4]
  assign _T_89507 = conflictPReg_9_9 ? 4'h9 : _T_89506; // @[LoadQueue.scala 191:60:@35933.4]
  assign _T_89508 = conflictPReg_9_10 ? 4'ha : _T_89507; // @[LoadQueue.scala 191:60:@35934.4]
  assign _T_89509 = conflictPReg_9_11 ? 4'hb : _T_89508; // @[LoadQueue.scala 191:60:@35935.4]
  assign _T_89510 = conflictPReg_9_12 ? 4'hc : _T_89509; // @[LoadQueue.scala 191:60:@35936.4]
  assign _T_89511 = conflictPReg_9_13 ? 4'hd : _T_89510; // @[LoadQueue.scala 191:60:@35937.4]
  assign _T_89512 = conflictPReg_9_14 ? 4'he : _T_89511; // @[LoadQueue.scala 191:60:@35938.4]
  assign _T_89513 = conflictPReg_9_15 ? 4'hf : _T_89512; // @[LoadQueue.scala 191:60:@35939.4]
  assign _T_89516 = conflictPReg_9_0 | conflictPReg_9_1; // @[LoadQueue.scala 192:43:@35941.4]
  assign _T_89517 = _T_89516 | conflictPReg_9_2; // @[LoadQueue.scala 192:43:@35942.4]
  assign _T_89518 = _T_89517 | conflictPReg_9_3; // @[LoadQueue.scala 192:43:@35943.4]
  assign _T_89519 = _T_89518 | conflictPReg_9_4; // @[LoadQueue.scala 192:43:@35944.4]
  assign _T_89520 = _T_89519 | conflictPReg_9_5; // @[LoadQueue.scala 192:43:@35945.4]
  assign _T_89521 = _T_89520 | conflictPReg_9_6; // @[LoadQueue.scala 192:43:@35946.4]
  assign _T_89522 = _T_89521 | conflictPReg_9_7; // @[LoadQueue.scala 192:43:@35947.4]
  assign _T_89523 = _T_89522 | conflictPReg_9_8; // @[LoadQueue.scala 192:43:@35948.4]
  assign _T_89524 = _T_89523 | conflictPReg_9_9; // @[LoadQueue.scala 192:43:@35949.4]
  assign _T_89525 = _T_89524 | conflictPReg_9_10; // @[LoadQueue.scala 192:43:@35950.4]
  assign _T_89526 = _T_89525 | conflictPReg_9_11; // @[LoadQueue.scala 192:43:@35951.4]
  assign _T_89527 = _T_89526 | conflictPReg_9_12; // @[LoadQueue.scala 192:43:@35952.4]
  assign _T_89528 = _T_89527 | conflictPReg_9_13; // @[LoadQueue.scala 192:43:@35953.4]
  assign _T_89529 = _T_89528 | conflictPReg_9_14; // @[LoadQueue.scala 192:43:@35954.4]
  assign _T_89530 = _T_89529 | conflictPReg_9_15; // @[LoadQueue.scala 192:43:@35955.4]
  assign _GEN_1458 = 4'h0 == _T_89513; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1459 = 4'h1 == _T_89513; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1460 = 4'h2 == _T_89513; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1461 = 4'h3 == _T_89513; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1462 = 4'h4 == _T_89513; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1463 = 4'h5 == _T_89513; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1464 = 4'h6 == _T_89513; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1465 = 4'h7 == _T_89513; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1466 = 4'h8 == _T_89513; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1467 = 4'h9 == _T_89513; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1468 = 4'ha == _T_89513; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1469 = 4'hb == _T_89513; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1470 = 4'hc == _T_89513; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1471 = 4'hd == _T_89513; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1472 = 4'he == _T_89513; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1473 = 4'hf == _T_89513; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1475 = 4'h1 == _T_89513 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1476 = 4'h2 == _T_89513 ? shiftedStoreDataKnownPReg_2 : _GEN_1475; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1477 = 4'h3 == _T_89513 ? shiftedStoreDataKnownPReg_3 : _GEN_1476; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1478 = 4'h4 == _T_89513 ? shiftedStoreDataKnownPReg_4 : _GEN_1477; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1479 = 4'h5 == _T_89513 ? shiftedStoreDataKnownPReg_5 : _GEN_1478; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1480 = 4'h6 == _T_89513 ? shiftedStoreDataKnownPReg_6 : _GEN_1479; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1481 = 4'h7 == _T_89513 ? shiftedStoreDataKnownPReg_7 : _GEN_1480; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1482 = 4'h8 == _T_89513 ? shiftedStoreDataKnownPReg_8 : _GEN_1481; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1483 = 4'h9 == _T_89513 ? shiftedStoreDataKnownPReg_9 : _GEN_1482; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1484 = 4'ha == _T_89513 ? shiftedStoreDataKnownPReg_10 : _GEN_1483; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1485 = 4'hb == _T_89513 ? shiftedStoreDataKnownPReg_11 : _GEN_1484; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1486 = 4'hc == _T_89513 ? shiftedStoreDataKnownPReg_12 : _GEN_1485; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1487 = 4'hd == _T_89513 ? shiftedStoreDataKnownPReg_13 : _GEN_1486; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1488 = 4'he == _T_89513 ? shiftedStoreDataKnownPReg_14 : _GEN_1487; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1489 = 4'hf == _T_89513 ? shiftedStoreDataKnownPReg_15 : _GEN_1488; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1491 = 4'h1 == _T_89513 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1492 = 4'h2 == _T_89513 ? shiftedStoreDataQPreg_2 : _GEN_1491; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1493 = 4'h3 == _T_89513 ? shiftedStoreDataQPreg_3 : _GEN_1492; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1494 = 4'h4 == _T_89513 ? shiftedStoreDataQPreg_4 : _GEN_1493; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1495 = 4'h5 == _T_89513 ? shiftedStoreDataQPreg_5 : _GEN_1494; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1496 = 4'h6 == _T_89513 ? shiftedStoreDataQPreg_6 : _GEN_1495; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1497 = 4'h7 == _T_89513 ? shiftedStoreDataQPreg_7 : _GEN_1496; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1498 = 4'h8 == _T_89513 ? shiftedStoreDataQPreg_8 : _GEN_1497; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1499 = 4'h9 == _T_89513 ? shiftedStoreDataQPreg_9 : _GEN_1498; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1500 = 4'ha == _T_89513 ? shiftedStoreDataQPreg_10 : _GEN_1499; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1501 = 4'hb == _T_89513 ? shiftedStoreDataQPreg_11 : _GEN_1500; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1502 = 4'hc == _T_89513 ? shiftedStoreDataQPreg_12 : _GEN_1501; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1503 = 4'hd == _T_89513 ? shiftedStoreDataQPreg_13 : _GEN_1502; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1504 = 4'he == _T_89513 ? shiftedStoreDataQPreg_14 : _GEN_1503; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1505 = 4'hf == _T_89513 ? shiftedStoreDataQPreg_15 : _GEN_1504; // @[LoadQueue.scala 195:31:@35959.6]
  assign lastConflict_9_0 = _T_89530 ? _GEN_1458 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_1 = _T_89530 ? _GEN_1459 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_2 = _T_89530 ? _GEN_1460 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_3 = _T_89530 ? _GEN_1461 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_4 = _T_89530 ? _GEN_1462 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_5 = _T_89530 ? _GEN_1463 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_6 = _T_89530 ? _GEN_1464 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_7 = _T_89530 ? _GEN_1465 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_8 = _T_89530 ? _GEN_1466 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_9 = _T_89530 ? _GEN_1467 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_10 = _T_89530 ? _GEN_1468 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_11 = _T_89530 ? _GEN_1469 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_12 = _T_89530 ? _GEN_1470 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_13 = _T_89530 ? _GEN_1471 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_14 = _T_89530 ? _GEN_1472 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_15 = _T_89530 ? _GEN_1473 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign canBypass_9 = _T_89530 ? _GEN_1489 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign bypassVal_9 = _T_89530 ? _GEN_1505 : 32'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign _T_89636 = conflictPReg_10_2 ? 2'h2 : {{1'd0}, conflictPReg_10_1}; // @[LoadQueue.scala 191:60:@36013.4]
  assign _T_89637 = conflictPReg_10_3 ? 2'h3 : _T_89636; // @[LoadQueue.scala 191:60:@36014.4]
  assign _T_89638 = conflictPReg_10_4 ? 3'h4 : {{1'd0}, _T_89637}; // @[LoadQueue.scala 191:60:@36015.4]
  assign _T_89639 = conflictPReg_10_5 ? 3'h5 : _T_89638; // @[LoadQueue.scala 191:60:@36016.4]
  assign _T_89640 = conflictPReg_10_6 ? 3'h6 : _T_89639; // @[LoadQueue.scala 191:60:@36017.4]
  assign _T_89641 = conflictPReg_10_7 ? 3'h7 : _T_89640; // @[LoadQueue.scala 191:60:@36018.4]
  assign _T_89642 = conflictPReg_10_8 ? 4'h8 : {{1'd0}, _T_89641}; // @[LoadQueue.scala 191:60:@36019.4]
  assign _T_89643 = conflictPReg_10_9 ? 4'h9 : _T_89642; // @[LoadQueue.scala 191:60:@36020.4]
  assign _T_89644 = conflictPReg_10_10 ? 4'ha : _T_89643; // @[LoadQueue.scala 191:60:@36021.4]
  assign _T_89645 = conflictPReg_10_11 ? 4'hb : _T_89644; // @[LoadQueue.scala 191:60:@36022.4]
  assign _T_89646 = conflictPReg_10_12 ? 4'hc : _T_89645; // @[LoadQueue.scala 191:60:@36023.4]
  assign _T_89647 = conflictPReg_10_13 ? 4'hd : _T_89646; // @[LoadQueue.scala 191:60:@36024.4]
  assign _T_89648 = conflictPReg_10_14 ? 4'he : _T_89647; // @[LoadQueue.scala 191:60:@36025.4]
  assign _T_89649 = conflictPReg_10_15 ? 4'hf : _T_89648; // @[LoadQueue.scala 191:60:@36026.4]
  assign _T_89652 = conflictPReg_10_0 | conflictPReg_10_1; // @[LoadQueue.scala 192:43:@36028.4]
  assign _T_89653 = _T_89652 | conflictPReg_10_2; // @[LoadQueue.scala 192:43:@36029.4]
  assign _T_89654 = _T_89653 | conflictPReg_10_3; // @[LoadQueue.scala 192:43:@36030.4]
  assign _T_89655 = _T_89654 | conflictPReg_10_4; // @[LoadQueue.scala 192:43:@36031.4]
  assign _T_89656 = _T_89655 | conflictPReg_10_5; // @[LoadQueue.scala 192:43:@36032.4]
  assign _T_89657 = _T_89656 | conflictPReg_10_6; // @[LoadQueue.scala 192:43:@36033.4]
  assign _T_89658 = _T_89657 | conflictPReg_10_7; // @[LoadQueue.scala 192:43:@36034.4]
  assign _T_89659 = _T_89658 | conflictPReg_10_8; // @[LoadQueue.scala 192:43:@36035.4]
  assign _T_89660 = _T_89659 | conflictPReg_10_9; // @[LoadQueue.scala 192:43:@36036.4]
  assign _T_89661 = _T_89660 | conflictPReg_10_10; // @[LoadQueue.scala 192:43:@36037.4]
  assign _T_89662 = _T_89661 | conflictPReg_10_11; // @[LoadQueue.scala 192:43:@36038.4]
  assign _T_89663 = _T_89662 | conflictPReg_10_12; // @[LoadQueue.scala 192:43:@36039.4]
  assign _T_89664 = _T_89663 | conflictPReg_10_13; // @[LoadQueue.scala 192:43:@36040.4]
  assign _T_89665 = _T_89664 | conflictPReg_10_14; // @[LoadQueue.scala 192:43:@36041.4]
  assign _T_89666 = _T_89665 | conflictPReg_10_15; // @[LoadQueue.scala 192:43:@36042.4]
  assign _GEN_1524 = 4'h0 == _T_89649; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1525 = 4'h1 == _T_89649; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1526 = 4'h2 == _T_89649; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1527 = 4'h3 == _T_89649; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1528 = 4'h4 == _T_89649; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1529 = 4'h5 == _T_89649; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1530 = 4'h6 == _T_89649; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1531 = 4'h7 == _T_89649; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1532 = 4'h8 == _T_89649; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1533 = 4'h9 == _T_89649; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1534 = 4'ha == _T_89649; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1535 = 4'hb == _T_89649; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1536 = 4'hc == _T_89649; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1537 = 4'hd == _T_89649; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1538 = 4'he == _T_89649; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1539 = 4'hf == _T_89649; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1541 = 4'h1 == _T_89649 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1542 = 4'h2 == _T_89649 ? shiftedStoreDataKnownPReg_2 : _GEN_1541; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1543 = 4'h3 == _T_89649 ? shiftedStoreDataKnownPReg_3 : _GEN_1542; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1544 = 4'h4 == _T_89649 ? shiftedStoreDataKnownPReg_4 : _GEN_1543; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1545 = 4'h5 == _T_89649 ? shiftedStoreDataKnownPReg_5 : _GEN_1544; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1546 = 4'h6 == _T_89649 ? shiftedStoreDataKnownPReg_6 : _GEN_1545; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1547 = 4'h7 == _T_89649 ? shiftedStoreDataKnownPReg_7 : _GEN_1546; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1548 = 4'h8 == _T_89649 ? shiftedStoreDataKnownPReg_8 : _GEN_1547; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1549 = 4'h9 == _T_89649 ? shiftedStoreDataKnownPReg_9 : _GEN_1548; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1550 = 4'ha == _T_89649 ? shiftedStoreDataKnownPReg_10 : _GEN_1549; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1551 = 4'hb == _T_89649 ? shiftedStoreDataKnownPReg_11 : _GEN_1550; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1552 = 4'hc == _T_89649 ? shiftedStoreDataKnownPReg_12 : _GEN_1551; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1553 = 4'hd == _T_89649 ? shiftedStoreDataKnownPReg_13 : _GEN_1552; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1554 = 4'he == _T_89649 ? shiftedStoreDataKnownPReg_14 : _GEN_1553; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1555 = 4'hf == _T_89649 ? shiftedStoreDataKnownPReg_15 : _GEN_1554; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1557 = 4'h1 == _T_89649 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1558 = 4'h2 == _T_89649 ? shiftedStoreDataQPreg_2 : _GEN_1557; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1559 = 4'h3 == _T_89649 ? shiftedStoreDataQPreg_3 : _GEN_1558; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1560 = 4'h4 == _T_89649 ? shiftedStoreDataQPreg_4 : _GEN_1559; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1561 = 4'h5 == _T_89649 ? shiftedStoreDataQPreg_5 : _GEN_1560; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1562 = 4'h6 == _T_89649 ? shiftedStoreDataQPreg_6 : _GEN_1561; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1563 = 4'h7 == _T_89649 ? shiftedStoreDataQPreg_7 : _GEN_1562; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1564 = 4'h8 == _T_89649 ? shiftedStoreDataQPreg_8 : _GEN_1563; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1565 = 4'h9 == _T_89649 ? shiftedStoreDataQPreg_9 : _GEN_1564; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1566 = 4'ha == _T_89649 ? shiftedStoreDataQPreg_10 : _GEN_1565; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1567 = 4'hb == _T_89649 ? shiftedStoreDataQPreg_11 : _GEN_1566; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1568 = 4'hc == _T_89649 ? shiftedStoreDataQPreg_12 : _GEN_1567; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1569 = 4'hd == _T_89649 ? shiftedStoreDataQPreg_13 : _GEN_1568; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1570 = 4'he == _T_89649 ? shiftedStoreDataQPreg_14 : _GEN_1569; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1571 = 4'hf == _T_89649 ? shiftedStoreDataQPreg_15 : _GEN_1570; // @[LoadQueue.scala 195:31:@36046.6]
  assign lastConflict_10_0 = _T_89666 ? _GEN_1524 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_1 = _T_89666 ? _GEN_1525 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_2 = _T_89666 ? _GEN_1526 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_3 = _T_89666 ? _GEN_1527 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_4 = _T_89666 ? _GEN_1528 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_5 = _T_89666 ? _GEN_1529 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_6 = _T_89666 ? _GEN_1530 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_7 = _T_89666 ? _GEN_1531 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_8 = _T_89666 ? _GEN_1532 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_9 = _T_89666 ? _GEN_1533 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_10 = _T_89666 ? _GEN_1534 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_11 = _T_89666 ? _GEN_1535 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_12 = _T_89666 ? _GEN_1536 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_13 = _T_89666 ? _GEN_1537 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_14 = _T_89666 ? _GEN_1538 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_15 = _T_89666 ? _GEN_1539 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign canBypass_10 = _T_89666 ? _GEN_1555 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign bypassVal_10 = _T_89666 ? _GEN_1571 : 32'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign _T_89772 = conflictPReg_11_2 ? 2'h2 : {{1'd0}, conflictPReg_11_1}; // @[LoadQueue.scala 191:60:@36100.4]
  assign _T_89773 = conflictPReg_11_3 ? 2'h3 : _T_89772; // @[LoadQueue.scala 191:60:@36101.4]
  assign _T_89774 = conflictPReg_11_4 ? 3'h4 : {{1'd0}, _T_89773}; // @[LoadQueue.scala 191:60:@36102.4]
  assign _T_89775 = conflictPReg_11_5 ? 3'h5 : _T_89774; // @[LoadQueue.scala 191:60:@36103.4]
  assign _T_89776 = conflictPReg_11_6 ? 3'h6 : _T_89775; // @[LoadQueue.scala 191:60:@36104.4]
  assign _T_89777 = conflictPReg_11_7 ? 3'h7 : _T_89776; // @[LoadQueue.scala 191:60:@36105.4]
  assign _T_89778 = conflictPReg_11_8 ? 4'h8 : {{1'd0}, _T_89777}; // @[LoadQueue.scala 191:60:@36106.4]
  assign _T_89779 = conflictPReg_11_9 ? 4'h9 : _T_89778; // @[LoadQueue.scala 191:60:@36107.4]
  assign _T_89780 = conflictPReg_11_10 ? 4'ha : _T_89779; // @[LoadQueue.scala 191:60:@36108.4]
  assign _T_89781 = conflictPReg_11_11 ? 4'hb : _T_89780; // @[LoadQueue.scala 191:60:@36109.4]
  assign _T_89782 = conflictPReg_11_12 ? 4'hc : _T_89781; // @[LoadQueue.scala 191:60:@36110.4]
  assign _T_89783 = conflictPReg_11_13 ? 4'hd : _T_89782; // @[LoadQueue.scala 191:60:@36111.4]
  assign _T_89784 = conflictPReg_11_14 ? 4'he : _T_89783; // @[LoadQueue.scala 191:60:@36112.4]
  assign _T_89785 = conflictPReg_11_15 ? 4'hf : _T_89784; // @[LoadQueue.scala 191:60:@36113.4]
  assign _T_89788 = conflictPReg_11_0 | conflictPReg_11_1; // @[LoadQueue.scala 192:43:@36115.4]
  assign _T_89789 = _T_89788 | conflictPReg_11_2; // @[LoadQueue.scala 192:43:@36116.4]
  assign _T_89790 = _T_89789 | conflictPReg_11_3; // @[LoadQueue.scala 192:43:@36117.4]
  assign _T_89791 = _T_89790 | conflictPReg_11_4; // @[LoadQueue.scala 192:43:@36118.4]
  assign _T_89792 = _T_89791 | conflictPReg_11_5; // @[LoadQueue.scala 192:43:@36119.4]
  assign _T_89793 = _T_89792 | conflictPReg_11_6; // @[LoadQueue.scala 192:43:@36120.4]
  assign _T_89794 = _T_89793 | conflictPReg_11_7; // @[LoadQueue.scala 192:43:@36121.4]
  assign _T_89795 = _T_89794 | conflictPReg_11_8; // @[LoadQueue.scala 192:43:@36122.4]
  assign _T_89796 = _T_89795 | conflictPReg_11_9; // @[LoadQueue.scala 192:43:@36123.4]
  assign _T_89797 = _T_89796 | conflictPReg_11_10; // @[LoadQueue.scala 192:43:@36124.4]
  assign _T_89798 = _T_89797 | conflictPReg_11_11; // @[LoadQueue.scala 192:43:@36125.4]
  assign _T_89799 = _T_89798 | conflictPReg_11_12; // @[LoadQueue.scala 192:43:@36126.4]
  assign _T_89800 = _T_89799 | conflictPReg_11_13; // @[LoadQueue.scala 192:43:@36127.4]
  assign _T_89801 = _T_89800 | conflictPReg_11_14; // @[LoadQueue.scala 192:43:@36128.4]
  assign _T_89802 = _T_89801 | conflictPReg_11_15; // @[LoadQueue.scala 192:43:@36129.4]
  assign _GEN_1590 = 4'h0 == _T_89785; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1591 = 4'h1 == _T_89785; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1592 = 4'h2 == _T_89785; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1593 = 4'h3 == _T_89785; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1594 = 4'h4 == _T_89785; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1595 = 4'h5 == _T_89785; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1596 = 4'h6 == _T_89785; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1597 = 4'h7 == _T_89785; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1598 = 4'h8 == _T_89785; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1599 = 4'h9 == _T_89785; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1600 = 4'ha == _T_89785; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1601 = 4'hb == _T_89785; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1602 = 4'hc == _T_89785; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1603 = 4'hd == _T_89785; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1604 = 4'he == _T_89785; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1605 = 4'hf == _T_89785; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1607 = 4'h1 == _T_89785 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1608 = 4'h2 == _T_89785 ? shiftedStoreDataKnownPReg_2 : _GEN_1607; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1609 = 4'h3 == _T_89785 ? shiftedStoreDataKnownPReg_3 : _GEN_1608; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1610 = 4'h4 == _T_89785 ? shiftedStoreDataKnownPReg_4 : _GEN_1609; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1611 = 4'h5 == _T_89785 ? shiftedStoreDataKnownPReg_5 : _GEN_1610; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1612 = 4'h6 == _T_89785 ? shiftedStoreDataKnownPReg_6 : _GEN_1611; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1613 = 4'h7 == _T_89785 ? shiftedStoreDataKnownPReg_7 : _GEN_1612; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1614 = 4'h8 == _T_89785 ? shiftedStoreDataKnownPReg_8 : _GEN_1613; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1615 = 4'h9 == _T_89785 ? shiftedStoreDataKnownPReg_9 : _GEN_1614; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1616 = 4'ha == _T_89785 ? shiftedStoreDataKnownPReg_10 : _GEN_1615; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1617 = 4'hb == _T_89785 ? shiftedStoreDataKnownPReg_11 : _GEN_1616; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1618 = 4'hc == _T_89785 ? shiftedStoreDataKnownPReg_12 : _GEN_1617; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1619 = 4'hd == _T_89785 ? shiftedStoreDataKnownPReg_13 : _GEN_1618; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1620 = 4'he == _T_89785 ? shiftedStoreDataKnownPReg_14 : _GEN_1619; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1621 = 4'hf == _T_89785 ? shiftedStoreDataKnownPReg_15 : _GEN_1620; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1623 = 4'h1 == _T_89785 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1624 = 4'h2 == _T_89785 ? shiftedStoreDataQPreg_2 : _GEN_1623; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1625 = 4'h3 == _T_89785 ? shiftedStoreDataQPreg_3 : _GEN_1624; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1626 = 4'h4 == _T_89785 ? shiftedStoreDataQPreg_4 : _GEN_1625; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1627 = 4'h5 == _T_89785 ? shiftedStoreDataQPreg_5 : _GEN_1626; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1628 = 4'h6 == _T_89785 ? shiftedStoreDataQPreg_6 : _GEN_1627; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1629 = 4'h7 == _T_89785 ? shiftedStoreDataQPreg_7 : _GEN_1628; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1630 = 4'h8 == _T_89785 ? shiftedStoreDataQPreg_8 : _GEN_1629; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1631 = 4'h9 == _T_89785 ? shiftedStoreDataQPreg_9 : _GEN_1630; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1632 = 4'ha == _T_89785 ? shiftedStoreDataQPreg_10 : _GEN_1631; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1633 = 4'hb == _T_89785 ? shiftedStoreDataQPreg_11 : _GEN_1632; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1634 = 4'hc == _T_89785 ? shiftedStoreDataQPreg_12 : _GEN_1633; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1635 = 4'hd == _T_89785 ? shiftedStoreDataQPreg_13 : _GEN_1634; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1636 = 4'he == _T_89785 ? shiftedStoreDataQPreg_14 : _GEN_1635; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1637 = 4'hf == _T_89785 ? shiftedStoreDataQPreg_15 : _GEN_1636; // @[LoadQueue.scala 195:31:@36133.6]
  assign lastConflict_11_0 = _T_89802 ? _GEN_1590 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_1 = _T_89802 ? _GEN_1591 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_2 = _T_89802 ? _GEN_1592 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_3 = _T_89802 ? _GEN_1593 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_4 = _T_89802 ? _GEN_1594 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_5 = _T_89802 ? _GEN_1595 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_6 = _T_89802 ? _GEN_1596 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_7 = _T_89802 ? _GEN_1597 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_8 = _T_89802 ? _GEN_1598 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_9 = _T_89802 ? _GEN_1599 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_10 = _T_89802 ? _GEN_1600 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_11 = _T_89802 ? _GEN_1601 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_12 = _T_89802 ? _GEN_1602 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_13 = _T_89802 ? _GEN_1603 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_14 = _T_89802 ? _GEN_1604 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_15 = _T_89802 ? _GEN_1605 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign canBypass_11 = _T_89802 ? _GEN_1621 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign bypassVal_11 = _T_89802 ? _GEN_1637 : 32'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign _T_89908 = conflictPReg_12_2 ? 2'h2 : {{1'd0}, conflictPReg_12_1}; // @[LoadQueue.scala 191:60:@36187.4]
  assign _T_89909 = conflictPReg_12_3 ? 2'h3 : _T_89908; // @[LoadQueue.scala 191:60:@36188.4]
  assign _T_89910 = conflictPReg_12_4 ? 3'h4 : {{1'd0}, _T_89909}; // @[LoadQueue.scala 191:60:@36189.4]
  assign _T_89911 = conflictPReg_12_5 ? 3'h5 : _T_89910; // @[LoadQueue.scala 191:60:@36190.4]
  assign _T_89912 = conflictPReg_12_6 ? 3'h6 : _T_89911; // @[LoadQueue.scala 191:60:@36191.4]
  assign _T_89913 = conflictPReg_12_7 ? 3'h7 : _T_89912; // @[LoadQueue.scala 191:60:@36192.4]
  assign _T_89914 = conflictPReg_12_8 ? 4'h8 : {{1'd0}, _T_89913}; // @[LoadQueue.scala 191:60:@36193.4]
  assign _T_89915 = conflictPReg_12_9 ? 4'h9 : _T_89914; // @[LoadQueue.scala 191:60:@36194.4]
  assign _T_89916 = conflictPReg_12_10 ? 4'ha : _T_89915; // @[LoadQueue.scala 191:60:@36195.4]
  assign _T_89917 = conflictPReg_12_11 ? 4'hb : _T_89916; // @[LoadQueue.scala 191:60:@36196.4]
  assign _T_89918 = conflictPReg_12_12 ? 4'hc : _T_89917; // @[LoadQueue.scala 191:60:@36197.4]
  assign _T_89919 = conflictPReg_12_13 ? 4'hd : _T_89918; // @[LoadQueue.scala 191:60:@36198.4]
  assign _T_89920 = conflictPReg_12_14 ? 4'he : _T_89919; // @[LoadQueue.scala 191:60:@36199.4]
  assign _T_89921 = conflictPReg_12_15 ? 4'hf : _T_89920; // @[LoadQueue.scala 191:60:@36200.4]
  assign _T_89924 = conflictPReg_12_0 | conflictPReg_12_1; // @[LoadQueue.scala 192:43:@36202.4]
  assign _T_89925 = _T_89924 | conflictPReg_12_2; // @[LoadQueue.scala 192:43:@36203.4]
  assign _T_89926 = _T_89925 | conflictPReg_12_3; // @[LoadQueue.scala 192:43:@36204.4]
  assign _T_89927 = _T_89926 | conflictPReg_12_4; // @[LoadQueue.scala 192:43:@36205.4]
  assign _T_89928 = _T_89927 | conflictPReg_12_5; // @[LoadQueue.scala 192:43:@36206.4]
  assign _T_89929 = _T_89928 | conflictPReg_12_6; // @[LoadQueue.scala 192:43:@36207.4]
  assign _T_89930 = _T_89929 | conflictPReg_12_7; // @[LoadQueue.scala 192:43:@36208.4]
  assign _T_89931 = _T_89930 | conflictPReg_12_8; // @[LoadQueue.scala 192:43:@36209.4]
  assign _T_89932 = _T_89931 | conflictPReg_12_9; // @[LoadQueue.scala 192:43:@36210.4]
  assign _T_89933 = _T_89932 | conflictPReg_12_10; // @[LoadQueue.scala 192:43:@36211.4]
  assign _T_89934 = _T_89933 | conflictPReg_12_11; // @[LoadQueue.scala 192:43:@36212.4]
  assign _T_89935 = _T_89934 | conflictPReg_12_12; // @[LoadQueue.scala 192:43:@36213.4]
  assign _T_89936 = _T_89935 | conflictPReg_12_13; // @[LoadQueue.scala 192:43:@36214.4]
  assign _T_89937 = _T_89936 | conflictPReg_12_14; // @[LoadQueue.scala 192:43:@36215.4]
  assign _T_89938 = _T_89937 | conflictPReg_12_15; // @[LoadQueue.scala 192:43:@36216.4]
  assign _GEN_1656 = 4'h0 == _T_89921; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1657 = 4'h1 == _T_89921; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1658 = 4'h2 == _T_89921; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1659 = 4'h3 == _T_89921; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1660 = 4'h4 == _T_89921; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1661 = 4'h5 == _T_89921; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1662 = 4'h6 == _T_89921; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1663 = 4'h7 == _T_89921; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1664 = 4'h8 == _T_89921; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1665 = 4'h9 == _T_89921; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1666 = 4'ha == _T_89921; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1667 = 4'hb == _T_89921; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1668 = 4'hc == _T_89921; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1669 = 4'hd == _T_89921; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1670 = 4'he == _T_89921; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1671 = 4'hf == _T_89921; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1673 = 4'h1 == _T_89921 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1674 = 4'h2 == _T_89921 ? shiftedStoreDataKnownPReg_2 : _GEN_1673; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1675 = 4'h3 == _T_89921 ? shiftedStoreDataKnownPReg_3 : _GEN_1674; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1676 = 4'h4 == _T_89921 ? shiftedStoreDataKnownPReg_4 : _GEN_1675; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1677 = 4'h5 == _T_89921 ? shiftedStoreDataKnownPReg_5 : _GEN_1676; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1678 = 4'h6 == _T_89921 ? shiftedStoreDataKnownPReg_6 : _GEN_1677; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1679 = 4'h7 == _T_89921 ? shiftedStoreDataKnownPReg_7 : _GEN_1678; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1680 = 4'h8 == _T_89921 ? shiftedStoreDataKnownPReg_8 : _GEN_1679; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1681 = 4'h9 == _T_89921 ? shiftedStoreDataKnownPReg_9 : _GEN_1680; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1682 = 4'ha == _T_89921 ? shiftedStoreDataKnownPReg_10 : _GEN_1681; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1683 = 4'hb == _T_89921 ? shiftedStoreDataKnownPReg_11 : _GEN_1682; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1684 = 4'hc == _T_89921 ? shiftedStoreDataKnownPReg_12 : _GEN_1683; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1685 = 4'hd == _T_89921 ? shiftedStoreDataKnownPReg_13 : _GEN_1684; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1686 = 4'he == _T_89921 ? shiftedStoreDataKnownPReg_14 : _GEN_1685; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1687 = 4'hf == _T_89921 ? shiftedStoreDataKnownPReg_15 : _GEN_1686; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1689 = 4'h1 == _T_89921 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1690 = 4'h2 == _T_89921 ? shiftedStoreDataQPreg_2 : _GEN_1689; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1691 = 4'h3 == _T_89921 ? shiftedStoreDataQPreg_3 : _GEN_1690; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1692 = 4'h4 == _T_89921 ? shiftedStoreDataQPreg_4 : _GEN_1691; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1693 = 4'h5 == _T_89921 ? shiftedStoreDataQPreg_5 : _GEN_1692; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1694 = 4'h6 == _T_89921 ? shiftedStoreDataQPreg_6 : _GEN_1693; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1695 = 4'h7 == _T_89921 ? shiftedStoreDataQPreg_7 : _GEN_1694; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1696 = 4'h8 == _T_89921 ? shiftedStoreDataQPreg_8 : _GEN_1695; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1697 = 4'h9 == _T_89921 ? shiftedStoreDataQPreg_9 : _GEN_1696; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1698 = 4'ha == _T_89921 ? shiftedStoreDataQPreg_10 : _GEN_1697; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1699 = 4'hb == _T_89921 ? shiftedStoreDataQPreg_11 : _GEN_1698; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1700 = 4'hc == _T_89921 ? shiftedStoreDataQPreg_12 : _GEN_1699; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1701 = 4'hd == _T_89921 ? shiftedStoreDataQPreg_13 : _GEN_1700; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1702 = 4'he == _T_89921 ? shiftedStoreDataQPreg_14 : _GEN_1701; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1703 = 4'hf == _T_89921 ? shiftedStoreDataQPreg_15 : _GEN_1702; // @[LoadQueue.scala 195:31:@36220.6]
  assign lastConflict_12_0 = _T_89938 ? _GEN_1656 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_1 = _T_89938 ? _GEN_1657 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_2 = _T_89938 ? _GEN_1658 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_3 = _T_89938 ? _GEN_1659 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_4 = _T_89938 ? _GEN_1660 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_5 = _T_89938 ? _GEN_1661 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_6 = _T_89938 ? _GEN_1662 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_7 = _T_89938 ? _GEN_1663 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_8 = _T_89938 ? _GEN_1664 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_9 = _T_89938 ? _GEN_1665 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_10 = _T_89938 ? _GEN_1666 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_11 = _T_89938 ? _GEN_1667 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_12 = _T_89938 ? _GEN_1668 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_13 = _T_89938 ? _GEN_1669 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_14 = _T_89938 ? _GEN_1670 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_15 = _T_89938 ? _GEN_1671 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign canBypass_12 = _T_89938 ? _GEN_1687 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign bypassVal_12 = _T_89938 ? _GEN_1703 : 32'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign _T_90044 = conflictPReg_13_2 ? 2'h2 : {{1'd0}, conflictPReg_13_1}; // @[LoadQueue.scala 191:60:@36274.4]
  assign _T_90045 = conflictPReg_13_3 ? 2'h3 : _T_90044; // @[LoadQueue.scala 191:60:@36275.4]
  assign _T_90046 = conflictPReg_13_4 ? 3'h4 : {{1'd0}, _T_90045}; // @[LoadQueue.scala 191:60:@36276.4]
  assign _T_90047 = conflictPReg_13_5 ? 3'h5 : _T_90046; // @[LoadQueue.scala 191:60:@36277.4]
  assign _T_90048 = conflictPReg_13_6 ? 3'h6 : _T_90047; // @[LoadQueue.scala 191:60:@36278.4]
  assign _T_90049 = conflictPReg_13_7 ? 3'h7 : _T_90048; // @[LoadQueue.scala 191:60:@36279.4]
  assign _T_90050 = conflictPReg_13_8 ? 4'h8 : {{1'd0}, _T_90049}; // @[LoadQueue.scala 191:60:@36280.4]
  assign _T_90051 = conflictPReg_13_9 ? 4'h9 : _T_90050; // @[LoadQueue.scala 191:60:@36281.4]
  assign _T_90052 = conflictPReg_13_10 ? 4'ha : _T_90051; // @[LoadQueue.scala 191:60:@36282.4]
  assign _T_90053 = conflictPReg_13_11 ? 4'hb : _T_90052; // @[LoadQueue.scala 191:60:@36283.4]
  assign _T_90054 = conflictPReg_13_12 ? 4'hc : _T_90053; // @[LoadQueue.scala 191:60:@36284.4]
  assign _T_90055 = conflictPReg_13_13 ? 4'hd : _T_90054; // @[LoadQueue.scala 191:60:@36285.4]
  assign _T_90056 = conflictPReg_13_14 ? 4'he : _T_90055; // @[LoadQueue.scala 191:60:@36286.4]
  assign _T_90057 = conflictPReg_13_15 ? 4'hf : _T_90056; // @[LoadQueue.scala 191:60:@36287.4]
  assign _T_90060 = conflictPReg_13_0 | conflictPReg_13_1; // @[LoadQueue.scala 192:43:@36289.4]
  assign _T_90061 = _T_90060 | conflictPReg_13_2; // @[LoadQueue.scala 192:43:@36290.4]
  assign _T_90062 = _T_90061 | conflictPReg_13_3; // @[LoadQueue.scala 192:43:@36291.4]
  assign _T_90063 = _T_90062 | conflictPReg_13_4; // @[LoadQueue.scala 192:43:@36292.4]
  assign _T_90064 = _T_90063 | conflictPReg_13_5; // @[LoadQueue.scala 192:43:@36293.4]
  assign _T_90065 = _T_90064 | conflictPReg_13_6; // @[LoadQueue.scala 192:43:@36294.4]
  assign _T_90066 = _T_90065 | conflictPReg_13_7; // @[LoadQueue.scala 192:43:@36295.4]
  assign _T_90067 = _T_90066 | conflictPReg_13_8; // @[LoadQueue.scala 192:43:@36296.4]
  assign _T_90068 = _T_90067 | conflictPReg_13_9; // @[LoadQueue.scala 192:43:@36297.4]
  assign _T_90069 = _T_90068 | conflictPReg_13_10; // @[LoadQueue.scala 192:43:@36298.4]
  assign _T_90070 = _T_90069 | conflictPReg_13_11; // @[LoadQueue.scala 192:43:@36299.4]
  assign _T_90071 = _T_90070 | conflictPReg_13_12; // @[LoadQueue.scala 192:43:@36300.4]
  assign _T_90072 = _T_90071 | conflictPReg_13_13; // @[LoadQueue.scala 192:43:@36301.4]
  assign _T_90073 = _T_90072 | conflictPReg_13_14; // @[LoadQueue.scala 192:43:@36302.4]
  assign _T_90074 = _T_90073 | conflictPReg_13_15; // @[LoadQueue.scala 192:43:@36303.4]
  assign _GEN_1722 = 4'h0 == _T_90057; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1723 = 4'h1 == _T_90057; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1724 = 4'h2 == _T_90057; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1725 = 4'h3 == _T_90057; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1726 = 4'h4 == _T_90057; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1727 = 4'h5 == _T_90057; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1728 = 4'h6 == _T_90057; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1729 = 4'h7 == _T_90057; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1730 = 4'h8 == _T_90057; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1731 = 4'h9 == _T_90057; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1732 = 4'ha == _T_90057; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1733 = 4'hb == _T_90057; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1734 = 4'hc == _T_90057; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1735 = 4'hd == _T_90057; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1736 = 4'he == _T_90057; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1737 = 4'hf == _T_90057; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1739 = 4'h1 == _T_90057 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1740 = 4'h2 == _T_90057 ? shiftedStoreDataKnownPReg_2 : _GEN_1739; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1741 = 4'h3 == _T_90057 ? shiftedStoreDataKnownPReg_3 : _GEN_1740; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1742 = 4'h4 == _T_90057 ? shiftedStoreDataKnownPReg_4 : _GEN_1741; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1743 = 4'h5 == _T_90057 ? shiftedStoreDataKnownPReg_5 : _GEN_1742; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1744 = 4'h6 == _T_90057 ? shiftedStoreDataKnownPReg_6 : _GEN_1743; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1745 = 4'h7 == _T_90057 ? shiftedStoreDataKnownPReg_7 : _GEN_1744; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1746 = 4'h8 == _T_90057 ? shiftedStoreDataKnownPReg_8 : _GEN_1745; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1747 = 4'h9 == _T_90057 ? shiftedStoreDataKnownPReg_9 : _GEN_1746; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1748 = 4'ha == _T_90057 ? shiftedStoreDataKnownPReg_10 : _GEN_1747; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1749 = 4'hb == _T_90057 ? shiftedStoreDataKnownPReg_11 : _GEN_1748; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1750 = 4'hc == _T_90057 ? shiftedStoreDataKnownPReg_12 : _GEN_1749; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1751 = 4'hd == _T_90057 ? shiftedStoreDataKnownPReg_13 : _GEN_1750; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1752 = 4'he == _T_90057 ? shiftedStoreDataKnownPReg_14 : _GEN_1751; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1753 = 4'hf == _T_90057 ? shiftedStoreDataKnownPReg_15 : _GEN_1752; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1755 = 4'h1 == _T_90057 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1756 = 4'h2 == _T_90057 ? shiftedStoreDataQPreg_2 : _GEN_1755; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1757 = 4'h3 == _T_90057 ? shiftedStoreDataQPreg_3 : _GEN_1756; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1758 = 4'h4 == _T_90057 ? shiftedStoreDataQPreg_4 : _GEN_1757; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1759 = 4'h5 == _T_90057 ? shiftedStoreDataQPreg_5 : _GEN_1758; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1760 = 4'h6 == _T_90057 ? shiftedStoreDataQPreg_6 : _GEN_1759; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1761 = 4'h7 == _T_90057 ? shiftedStoreDataQPreg_7 : _GEN_1760; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1762 = 4'h8 == _T_90057 ? shiftedStoreDataQPreg_8 : _GEN_1761; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1763 = 4'h9 == _T_90057 ? shiftedStoreDataQPreg_9 : _GEN_1762; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1764 = 4'ha == _T_90057 ? shiftedStoreDataQPreg_10 : _GEN_1763; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1765 = 4'hb == _T_90057 ? shiftedStoreDataQPreg_11 : _GEN_1764; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1766 = 4'hc == _T_90057 ? shiftedStoreDataQPreg_12 : _GEN_1765; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1767 = 4'hd == _T_90057 ? shiftedStoreDataQPreg_13 : _GEN_1766; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1768 = 4'he == _T_90057 ? shiftedStoreDataQPreg_14 : _GEN_1767; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1769 = 4'hf == _T_90057 ? shiftedStoreDataQPreg_15 : _GEN_1768; // @[LoadQueue.scala 195:31:@36307.6]
  assign lastConflict_13_0 = _T_90074 ? _GEN_1722 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_1 = _T_90074 ? _GEN_1723 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_2 = _T_90074 ? _GEN_1724 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_3 = _T_90074 ? _GEN_1725 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_4 = _T_90074 ? _GEN_1726 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_5 = _T_90074 ? _GEN_1727 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_6 = _T_90074 ? _GEN_1728 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_7 = _T_90074 ? _GEN_1729 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_8 = _T_90074 ? _GEN_1730 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_9 = _T_90074 ? _GEN_1731 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_10 = _T_90074 ? _GEN_1732 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_11 = _T_90074 ? _GEN_1733 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_12 = _T_90074 ? _GEN_1734 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_13 = _T_90074 ? _GEN_1735 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_14 = _T_90074 ? _GEN_1736 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_15 = _T_90074 ? _GEN_1737 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign canBypass_13 = _T_90074 ? _GEN_1753 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign bypassVal_13 = _T_90074 ? _GEN_1769 : 32'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign _T_90180 = conflictPReg_14_2 ? 2'h2 : {{1'd0}, conflictPReg_14_1}; // @[LoadQueue.scala 191:60:@36361.4]
  assign _T_90181 = conflictPReg_14_3 ? 2'h3 : _T_90180; // @[LoadQueue.scala 191:60:@36362.4]
  assign _T_90182 = conflictPReg_14_4 ? 3'h4 : {{1'd0}, _T_90181}; // @[LoadQueue.scala 191:60:@36363.4]
  assign _T_90183 = conflictPReg_14_5 ? 3'h5 : _T_90182; // @[LoadQueue.scala 191:60:@36364.4]
  assign _T_90184 = conflictPReg_14_6 ? 3'h6 : _T_90183; // @[LoadQueue.scala 191:60:@36365.4]
  assign _T_90185 = conflictPReg_14_7 ? 3'h7 : _T_90184; // @[LoadQueue.scala 191:60:@36366.4]
  assign _T_90186 = conflictPReg_14_8 ? 4'h8 : {{1'd0}, _T_90185}; // @[LoadQueue.scala 191:60:@36367.4]
  assign _T_90187 = conflictPReg_14_9 ? 4'h9 : _T_90186; // @[LoadQueue.scala 191:60:@36368.4]
  assign _T_90188 = conflictPReg_14_10 ? 4'ha : _T_90187; // @[LoadQueue.scala 191:60:@36369.4]
  assign _T_90189 = conflictPReg_14_11 ? 4'hb : _T_90188; // @[LoadQueue.scala 191:60:@36370.4]
  assign _T_90190 = conflictPReg_14_12 ? 4'hc : _T_90189; // @[LoadQueue.scala 191:60:@36371.4]
  assign _T_90191 = conflictPReg_14_13 ? 4'hd : _T_90190; // @[LoadQueue.scala 191:60:@36372.4]
  assign _T_90192 = conflictPReg_14_14 ? 4'he : _T_90191; // @[LoadQueue.scala 191:60:@36373.4]
  assign _T_90193 = conflictPReg_14_15 ? 4'hf : _T_90192; // @[LoadQueue.scala 191:60:@36374.4]
  assign _T_90196 = conflictPReg_14_0 | conflictPReg_14_1; // @[LoadQueue.scala 192:43:@36376.4]
  assign _T_90197 = _T_90196 | conflictPReg_14_2; // @[LoadQueue.scala 192:43:@36377.4]
  assign _T_90198 = _T_90197 | conflictPReg_14_3; // @[LoadQueue.scala 192:43:@36378.4]
  assign _T_90199 = _T_90198 | conflictPReg_14_4; // @[LoadQueue.scala 192:43:@36379.4]
  assign _T_90200 = _T_90199 | conflictPReg_14_5; // @[LoadQueue.scala 192:43:@36380.4]
  assign _T_90201 = _T_90200 | conflictPReg_14_6; // @[LoadQueue.scala 192:43:@36381.4]
  assign _T_90202 = _T_90201 | conflictPReg_14_7; // @[LoadQueue.scala 192:43:@36382.4]
  assign _T_90203 = _T_90202 | conflictPReg_14_8; // @[LoadQueue.scala 192:43:@36383.4]
  assign _T_90204 = _T_90203 | conflictPReg_14_9; // @[LoadQueue.scala 192:43:@36384.4]
  assign _T_90205 = _T_90204 | conflictPReg_14_10; // @[LoadQueue.scala 192:43:@36385.4]
  assign _T_90206 = _T_90205 | conflictPReg_14_11; // @[LoadQueue.scala 192:43:@36386.4]
  assign _T_90207 = _T_90206 | conflictPReg_14_12; // @[LoadQueue.scala 192:43:@36387.4]
  assign _T_90208 = _T_90207 | conflictPReg_14_13; // @[LoadQueue.scala 192:43:@36388.4]
  assign _T_90209 = _T_90208 | conflictPReg_14_14; // @[LoadQueue.scala 192:43:@36389.4]
  assign _T_90210 = _T_90209 | conflictPReg_14_15; // @[LoadQueue.scala 192:43:@36390.4]
  assign _GEN_1788 = 4'h0 == _T_90193; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1789 = 4'h1 == _T_90193; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1790 = 4'h2 == _T_90193; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1791 = 4'h3 == _T_90193; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1792 = 4'h4 == _T_90193; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1793 = 4'h5 == _T_90193; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1794 = 4'h6 == _T_90193; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1795 = 4'h7 == _T_90193; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1796 = 4'h8 == _T_90193; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1797 = 4'h9 == _T_90193; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1798 = 4'ha == _T_90193; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1799 = 4'hb == _T_90193; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1800 = 4'hc == _T_90193; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1801 = 4'hd == _T_90193; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1802 = 4'he == _T_90193; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1803 = 4'hf == _T_90193; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1805 = 4'h1 == _T_90193 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1806 = 4'h2 == _T_90193 ? shiftedStoreDataKnownPReg_2 : _GEN_1805; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1807 = 4'h3 == _T_90193 ? shiftedStoreDataKnownPReg_3 : _GEN_1806; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1808 = 4'h4 == _T_90193 ? shiftedStoreDataKnownPReg_4 : _GEN_1807; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1809 = 4'h5 == _T_90193 ? shiftedStoreDataKnownPReg_5 : _GEN_1808; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1810 = 4'h6 == _T_90193 ? shiftedStoreDataKnownPReg_6 : _GEN_1809; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1811 = 4'h7 == _T_90193 ? shiftedStoreDataKnownPReg_7 : _GEN_1810; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1812 = 4'h8 == _T_90193 ? shiftedStoreDataKnownPReg_8 : _GEN_1811; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1813 = 4'h9 == _T_90193 ? shiftedStoreDataKnownPReg_9 : _GEN_1812; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1814 = 4'ha == _T_90193 ? shiftedStoreDataKnownPReg_10 : _GEN_1813; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1815 = 4'hb == _T_90193 ? shiftedStoreDataKnownPReg_11 : _GEN_1814; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1816 = 4'hc == _T_90193 ? shiftedStoreDataKnownPReg_12 : _GEN_1815; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1817 = 4'hd == _T_90193 ? shiftedStoreDataKnownPReg_13 : _GEN_1816; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1818 = 4'he == _T_90193 ? shiftedStoreDataKnownPReg_14 : _GEN_1817; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1819 = 4'hf == _T_90193 ? shiftedStoreDataKnownPReg_15 : _GEN_1818; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1821 = 4'h1 == _T_90193 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1822 = 4'h2 == _T_90193 ? shiftedStoreDataQPreg_2 : _GEN_1821; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1823 = 4'h3 == _T_90193 ? shiftedStoreDataQPreg_3 : _GEN_1822; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1824 = 4'h4 == _T_90193 ? shiftedStoreDataQPreg_4 : _GEN_1823; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1825 = 4'h5 == _T_90193 ? shiftedStoreDataQPreg_5 : _GEN_1824; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1826 = 4'h6 == _T_90193 ? shiftedStoreDataQPreg_6 : _GEN_1825; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1827 = 4'h7 == _T_90193 ? shiftedStoreDataQPreg_7 : _GEN_1826; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1828 = 4'h8 == _T_90193 ? shiftedStoreDataQPreg_8 : _GEN_1827; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1829 = 4'h9 == _T_90193 ? shiftedStoreDataQPreg_9 : _GEN_1828; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1830 = 4'ha == _T_90193 ? shiftedStoreDataQPreg_10 : _GEN_1829; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1831 = 4'hb == _T_90193 ? shiftedStoreDataQPreg_11 : _GEN_1830; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1832 = 4'hc == _T_90193 ? shiftedStoreDataQPreg_12 : _GEN_1831; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1833 = 4'hd == _T_90193 ? shiftedStoreDataQPreg_13 : _GEN_1832; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1834 = 4'he == _T_90193 ? shiftedStoreDataQPreg_14 : _GEN_1833; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1835 = 4'hf == _T_90193 ? shiftedStoreDataQPreg_15 : _GEN_1834; // @[LoadQueue.scala 195:31:@36394.6]
  assign lastConflict_14_0 = _T_90210 ? _GEN_1788 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_1 = _T_90210 ? _GEN_1789 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_2 = _T_90210 ? _GEN_1790 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_3 = _T_90210 ? _GEN_1791 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_4 = _T_90210 ? _GEN_1792 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_5 = _T_90210 ? _GEN_1793 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_6 = _T_90210 ? _GEN_1794 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_7 = _T_90210 ? _GEN_1795 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_8 = _T_90210 ? _GEN_1796 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_9 = _T_90210 ? _GEN_1797 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_10 = _T_90210 ? _GEN_1798 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_11 = _T_90210 ? _GEN_1799 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_12 = _T_90210 ? _GEN_1800 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_13 = _T_90210 ? _GEN_1801 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_14 = _T_90210 ? _GEN_1802 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_15 = _T_90210 ? _GEN_1803 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign canBypass_14 = _T_90210 ? _GEN_1819 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign bypassVal_14 = _T_90210 ? _GEN_1835 : 32'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign _T_90316 = conflictPReg_15_2 ? 2'h2 : {{1'd0}, conflictPReg_15_1}; // @[LoadQueue.scala 191:60:@36448.4]
  assign _T_90317 = conflictPReg_15_3 ? 2'h3 : _T_90316; // @[LoadQueue.scala 191:60:@36449.4]
  assign _T_90318 = conflictPReg_15_4 ? 3'h4 : {{1'd0}, _T_90317}; // @[LoadQueue.scala 191:60:@36450.4]
  assign _T_90319 = conflictPReg_15_5 ? 3'h5 : _T_90318; // @[LoadQueue.scala 191:60:@36451.4]
  assign _T_90320 = conflictPReg_15_6 ? 3'h6 : _T_90319; // @[LoadQueue.scala 191:60:@36452.4]
  assign _T_90321 = conflictPReg_15_7 ? 3'h7 : _T_90320; // @[LoadQueue.scala 191:60:@36453.4]
  assign _T_90322 = conflictPReg_15_8 ? 4'h8 : {{1'd0}, _T_90321}; // @[LoadQueue.scala 191:60:@36454.4]
  assign _T_90323 = conflictPReg_15_9 ? 4'h9 : _T_90322; // @[LoadQueue.scala 191:60:@36455.4]
  assign _T_90324 = conflictPReg_15_10 ? 4'ha : _T_90323; // @[LoadQueue.scala 191:60:@36456.4]
  assign _T_90325 = conflictPReg_15_11 ? 4'hb : _T_90324; // @[LoadQueue.scala 191:60:@36457.4]
  assign _T_90326 = conflictPReg_15_12 ? 4'hc : _T_90325; // @[LoadQueue.scala 191:60:@36458.4]
  assign _T_90327 = conflictPReg_15_13 ? 4'hd : _T_90326; // @[LoadQueue.scala 191:60:@36459.4]
  assign _T_90328 = conflictPReg_15_14 ? 4'he : _T_90327; // @[LoadQueue.scala 191:60:@36460.4]
  assign _T_90329 = conflictPReg_15_15 ? 4'hf : _T_90328; // @[LoadQueue.scala 191:60:@36461.4]
  assign _T_90332 = conflictPReg_15_0 | conflictPReg_15_1; // @[LoadQueue.scala 192:43:@36463.4]
  assign _T_90333 = _T_90332 | conflictPReg_15_2; // @[LoadQueue.scala 192:43:@36464.4]
  assign _T_90334 = _T_90333 | conflictPReg_15_3; // @[LoadQueue.scala 192:43:@36465.4]
  assign _T_90335 = _T_90334 | conflictPReg_15_4; // @[LoadQueue.scala 192:43:@36466.4]
  assign _T_90336 = _T_90335 | conflictPReg_15_5; // @[LoadQueue.scala 192:43:@36467.4]
  assign _T_90337 = _T_90336 | conflictPReg_15_6; // @[LoadQueue.scala 192:43:@36468.4]
  assign _T_90338 = _T_90337 | conflictPReg_15_7; // @[LoadQueue.scala 192:43:@36469.4]
  assign _T_90339 = _T_90338 | conflictPReg_15_8; // @[LoadQueue.scala 192:43:@36470.4]
  assign _T_90340 = _T_90339 | conflictPReg_15_9; // @[LoadQueue.scala 192:43:@36471.4]
  assign _T_90341 = _T_90340 | conflictPReg_15_10; // @[LoadQueue.scala 192:43:@36472.4]
  assign _T_90342 = _T_90341 | conflictPReg_15_11; // @[LoadQueue.scala 192:43:@36473.4]
  assign _T_90343 = _T_90342 | conflictPReg_15_12; // @[LoadQueue.scala 192:43:@36474.4]
  assign _T_90344 = _T_90343 | conflictPReg_15_13; // @[LoadQueue.scala 192:43:@36475.4]
  assign _T_90345 = _T_90344 | conflictPReg_15_14; // @[LoadQueue.scala 192:43:@36476.4]
  assign _T_90346 = _T_90345 | conflictPReg_15_15; // @[LoadQueue.scala 192:43:@36477.4]
  assign _GEN_1854 = 4'h0 == _T_90329; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1855 = 4'h1 == _T_90329; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1856 = 4'h2 == _T_90329; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1857 = 4'h3 == _T_90329; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1858 = 4'h4 == _T_90329; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1859 = 4'h5 == _T_90329; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1860 = 4'h6 == _T_90329; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1861 = 4'h7 == _T_90329; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1862 = 4'h8 == _T_90329; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1863 = 4'h9 == _T_90329; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1864 = 4'ha == _T_90329; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1865 = 4'hb == _T_90329; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1866 = 4'hc == _T_90329; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1867 = 4'hd == _T_90329; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1868 = 4'he == _T_90329; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1869 = 4'hf == _T_90329; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1871 = 4'h1 == _T_90329 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1872 = 4'h2 == _T_90329 ? shiftedStoreDataKnownPReg_2 : _GEN_1871; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1873 = 4'h3 == _T_90329 ? shiftedStoreDataKnownPReg_3 : _GEN_1872; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1874 = 4'h4 == _T_90329 ? shiftedStoreDataKnownPReg_4 : _GEN_1873; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1875 = 4'h5 == _T_90329 ? shiftedStoreDataKnownPReg_5 : _GEN_1874; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1876 = 4'h6 == _T_90329 ? shiftedStoreDataKnownPReg_6 : _GEN_1875; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1877 = 4'h7 == _T_90329 ? shiftedStoreDataKnownPReg_7 : _GEN_1876; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1878 = 4'h8 == _T_90329 ? shiftedStoreDataKnownPReg_8 : _GEN_1877; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1879 = 4'h9 == _T_90329 ? shiftedStoreDataKnownPReg_9 : _GEN_1878; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1880 = 4'ha == _T_90329 ? shiftedStoreDataKnownPReg_10 : _GEN_1879; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1881 = 4'hb == _T_90329 ? shiftedStoreDataKnownPReg_11 : _GEN_1880; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1882 = 4'hc == _T_90329 ? shiftedStoreDataKnownPReg_12 : _GEN_1881; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1883 = 4'hd == _T_90329 ? shiftedStoreDataKnownPReg_13 : _GEN_1882; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1884 = 4'he == _T_90329 ? shiftedStoreDataKnownPReg_14 : _GEN_1883; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1885 = 4'hf == _T_90329 ? shiftedStoreDataKnownPReg_15 : _GEN_1884; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1887 = 4'h1 == _T_90329 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1888 = 4'h2 == _T_90329 ? shiftedStoreDataQPreg_2 : _GEN_1887; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1889 = 4'h3 == _T_90329 ? shiftedStoreDataQPreg_3 : _GEN_1888; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1890 = 4'h4 == _T_90329 ? shiftedStoreDataQPreg_4 : _GEN_1889; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1891 = 4'h5 == _T_90329 ? shiftedStoreDataQPreg_5 : _GEN_1890; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1892 = 4'h6 == _T_90329 ? shiftedStoreDataQPreg_6 : _GEN_1891; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1893 = 4'h7 == _T_90329 ? shiftedStoreDataQPreg_7 : _GEN_1892; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1894 = 4'h8 == _T_90329 ? shiftedStoreDataQPreg_8 : _GEN_1893; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1895 = 4'h9 == _T_90329 ? shiftedStoreDataQPreg_9 : _GEN_1894; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1896 = 4'ha == _T_90329 ? shiftedStoreDataQPreg_10 : _GEN_1895; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1897 = 4'hb == _T_90329 ? shiftedStoreDataQPreg_11 : _GEN_1896; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1898 = 4'hc == _T_90329 ? shiftedStoreDataQPreg_12 : _GEN_1897; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1899 = 4'hd == _T_90329 ? shiftedStoreDataQPreg_13 : _GEN_1898; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1900 = 4'he == _T_90329 ? shiftedStoreDataQPreg_14 : _GEN_1899; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1901 = 4'hf == _T_90329 ? shiftedStoreDataQPreg_15 : _GEN_1900; // @[LoadQueue.scala 195:31:@36481.6]
  assign lastConflict_15_0 = _T_90346 ? _GEN_1854 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_1 = _T_90346 ? _GEN_1855 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_2 = _T_90346 ? _GEN_1856 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_3 = _T_90346 ? _GEN_1857 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_4 = _T_90346 ? _GEN_1858 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_5 = _T_90346 ? _GEN_1859 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_6 = _T_90346 ? _GEN_1860 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_7 = _T_90346 ? _GEN_1861 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_8 = _T_90346 ? _GEN_1862 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_9 = _T_90346 ? _GEN_1863 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_10 = _T_90346 ? _GEN_1864 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_11 = _T_90346 ? _GEN_1865 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_12 = _T_90346 ? _GEN_1866 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_13 = _T_90346 ? _GEN_1867 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_14 = _T_90346 ? _GEN_1868 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_15 = _T_90346 ? _GEN_1869 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign canBypass_15 = _T_90346 ? _GEN_1885 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign bypassVal_15 = _T_90346 ? _GEN_1901 : 32'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign _T_90406 = 16'h1 << head; // @[OneHot.scala 52:12:@36486.4]
  assign _T_90408 = _T_90406[0]; // @[util.scala 33:60:@36488.4]
  assign _T_90409 = _T_90406[1]; // @[util.scala 33:60:@36489.4]
  assign _T_90410 = _T_90406[2]; // @[util.scala 33:60:@36490.4]
  assign _T_90411 = _T_90406[3]; // @[util.scala 33:60:@36491.4]
  assign _T_90412 = _T_90406[4]; // @[util.scala 33:60:@36492.4]
  assign _T_90413 = _T_90406[5]; // @[util.scala 33:60:@36493.4]
  assign _T_90414 = _T_90406[6]; // @[util.scala 33:60:@36494.4]
  assign _T_90415 = _T_90406[7]; // @[util.scala 33:60:@36495.4]
  assign _T_90416 = _T_90406[8]; // @[util.scala 33:60:@36496.4]
  assign _T_90417 = _T_90406[9]; // @[util.scala 33:60:@36497.4]
  assign _T_90418 = _T_90406[10]; // @[util.scala 33:60:@36498.4]
  assign _T_90419 = _T_90406[11]; // @[util.scala 33:60:@36499.4]
  assign _T_90420 = _T_90406[12]; // @[util.scala 33:60:@36500.4]
  assign _T_90421 = _T_90406[13]; // @[util.scala 33:60:@36501.4]
  assign _T_90422 = _T_90406[14]; // @[util.scala 33:60:@36502.4]
  assign _T_90423 = _T_90406[15]; // @[util.scala 33:60:@36503.4]
  assign _T_93520 = dataKnownPReg_15 == 1'h0; // @[LoadQueue.scala 229:41:@39026.4]
  assign _T_93521 = addrKnownPReg_15 & _T_93520; // @[LoadQueue.scala 229:38:@39027.4]
  assign _T_93523 = bypassInitiated_15 == 1'h0; // @[LoadQueue.scala 230:12:@39029.6]
  assign _T_93525 = prevPriorityRequest_15 == 1'h0; // @[LoadQueue.scala 230:46:@39030.6]
  assign _T_93526 = _T_93523 & _T_93525; // @[LoadQueue.scala 230:43:@39031.6]
  assign _T_93528 = dataKnown_15 == 1'h0; // @[LoadQueue.scala 230:84:@39032.6]
  assign _T_93529 = _T_93526 & _T_93528; // @[LoadQueue.scala 230:81:@39033.6]
  assign _T_93532 = storeAddrNotKnownFlagsPReg_15_0 | storeAddrNotKnownFlagsPReg_15_1; // @[LoadQueue.scala 233:86:@39036.8]
  assign _T_93533 = _T_93532 | storeAddrNotKnownFlagsPReg_15_2; // @[LoadQueue.scala 233:86:@39037.8]
  assign _T_93534 = _T_93533 | storeAddrNotKnownFlagsPReg_15_3; // @[LoadQueue.scala 233:86:@39038.8]
  assign _T_93535 = _T_93534 | storeAddrNotKnownFlagsPReg_15_4; // @[LoadQueue.scala 233:86:@39039.8]
  assign _T_93536 = _T_93535 | storeAddrNotKnownFlagsPReg_15_5; // @[LoadQueue.scala 233:86:@39040.8]
  assign _T_93537 = _T_93536 | storeAddrNotKnownFlagsPReg_15_6; // @[LoadQueue.scala 233:86:@39041.8]
  assign _T_93538 = _T_93537 | storeAddrNotKnownFlagsPReg_15_7; // @[LoadQueue.scala 233:86:@39042.8]
  assign _T_93539 = _T_93538 | storeAddrNotKnownFlagsPReg_15_8; // @[LoadQueue.scala 233:86:@39043.8]
  assign _T_93540 = _T_93539 | storeAddrNotKnownFlagsPReg_15_9; // @[LoadQueue.scala 233:86:@39044.8]
  assign _T_93541 = _T_93540 | storeAddrNotKnownFlagsPReg_15_10; // @[LoadQueue.scala 233:86:@39045.8]
  assign _T_93542 = _T_93541 | storeAddrNotKnownFlagsPReg_15_11; // @[LoadQueue.scala 233:86:@39046.8]
  assign _T_93543 = _T_93542 | storeAddrNotKnownFlagsPReg_15_12; // @[LoadQueue.scala 233:86:@39047.8]
  assign _T_93544 = _T_93543 | storeAddrNotKnownFlagsPReg_15_13; // @[LoadQueue.scala 233:86:@39048.8]
  assign _T_93545 = _T_93544 | storeAddrNotKnownFlagsPReg_15_14; // @[LoadQueue.scala 233:86:@39049.8]
  assign _T_93546 = _T_93545 | storeAddrNotKnownFlagsPReg_15_15; // @[LoadQueue.scala 233:86:@39050.8]
  assign _T_93548 = _T_93546 == 1'h0; // @[LoadQueue.scala 233:38:@39051.8]
  assign _T_93567 = _T_90346 == 1'h0; // @[LoadQueue.scala 234:11:@39068.8]
  assign _T_93568 = _T_93548 & _T_93567; // @[LoadQueue.scala 233:103:@39069.8]
  assign _GEN_2028 = _T_93529 ? _T_93568 : 1'h0; // @[LoadQueue.scala 230:110:@39034.6]
  assign loadRequest_15 = _T_93521 ? _GEN_2028 : 1'h0; // @[LoadQueue.scala 229:71:@39028.4]
  assign _T_90464 = loadRequest_15 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36521.4]
  assign _T_93436 = dataKnownPReg_14 == 1'h0; // @[LoadQueue.scala 229:41:@38944.4]
  assign _T_93437 = addrKnownPReg_14 & _T_93436; // @[LoadQueue.scala 229:38:@38945.4]
  assign _T_93439 = bypassInitiated_14 == 1'h0; // @[LoadQueue.scala 230:12:@38947.6]
  assign _T_93441 = prevPriorityRequest_14 == 1'h0; // @[LoadQueue.scala 230:46:@38948.6]
  assign _T_93442 = _T_93439 & _T_93441; // @[LoadQueue.scala 230:43:@38949.6]
  assign _T_93444 = dataKnown_14 == 1'h0; // @[LoadQueue.scala 230:84:@38950.6]
  assign _T_93445 = _T_93442 & _T_93444; // @[LoadQueue.scala 230:81:@38951.6]
  assign _T_93448 = storeAddrNotKnownFlagsPReg_14_0 | storeAddrNotKnownFlagsPReg_14_1; // @[LoadQueue.scala 233:86:@38954.8]
  assign _T_93449 = _T_93448 | storeAddrNotKnownFlagsPReg_14_2; // @[LoadQueue.scala 233:86:@38955.8]
  assign _T_93450 = _T_93449 | storeAddrNotKnownFlagsPReg_14_3; // @[LoadQueue.scala 233:86:@38956.8]
  assign _T_93451 = _T_93450 | storeAddrNotKnownFlagsPReg_14_4; // @[LoadQueue.scala 233:86:@38957.8]
  assign _T_93452 = _T_93451 | storeAddrNotKnownFlagsPReg_14_5; // @[LoadQueue.scala 233:86:@38958.8]
  assign _T_93453 = _T_93452 | storeAddrNotKnownFlagsPReg_14_6; // @[LoadQueue.scala 233:86:@38959.8]
  assign _T_93454 = _T_93453 | storeAddrNotKnownFlagsPReg_14_7; // @[LoadQueue.scala 233:86:@38960.8]
  assign _T_93455 = _T_93454 | storeAddrNotKnownFlagsPReg_14_8; // @[LoadQueue.scala 233:86:@38961.8]
  assign _T_93456 = _T_93455 | storeAddrNotKnownFlagsPReg_14_9; // @[LoadQueue.scala 233:86:@38962.8]
  assign _T_93457 = _T_93456 | storeAddrNotKnownFlagsPReg_14_10; // @[LoadQueue.scala 233:86:@38963.8]
  assign _T_93458 = _T_93457 | storeAddrNotKnownFlagsPReg_14_11; // @[LoadQueue.scala 233:86:@38964.8]
  assign _T_93459 = _T_93458 | storeAddrNotKnownFlagsPReg_14_12; // @[LoadQueue.scala 233:86:@38965.8]
  assign _T_93460 = _T_93459 | storeAddrNotKnownFlagsPReg_14_13; // @[LoadQueue.scala 233:86:@38966.8]
  assign _T_93461 = _T_93460 | storeAddrNotKnownFlagsPReg_14_14; // @[LoadQueue.scala 233:86:@38967.8]
  assign _T_93462 = _T_93461 | storeAddrNotKnownFlagsPReg_14_15; // @[LoadQueue.scala 233:86:@38968.8]
  assign _T_93464 = _T_93462 == 1'h0; // @[LoadQueue.scala 233:38:@38969.8]
  assign _T_93483 = _T_90210 == 1'h0; // @[LoadQueue.scala 234:11:@38986.8]
  assign _T_93484 = _T_93464 & _T_93483; // @[LoadQueue.scala 233:103:@38987.8]
  assign _GEN_2024 = _T_93445 ? _T_93484 : 1'h0; // @[LoadQueue.scala 230:110:@38952.6]
  assign loadRequest_14 = _T_93437 ? _GEN_2024 : 1'h0; // @[LoadQueue.scala 229:71:@38946.4]
  assign _T_90465 = loadRequest_14 ? 16'h4000 : _T_90464; // @[Mux.scala 31:69:@36522.4]
  assign _T_93352 = dataKnownPReg_13 == 1'h0; // @[LoadQueue.scala 229:41:@38862.4]
  assign _T_93353 = addrKnownPReg_13 & _T_93352; // @[LoadQueue.scala 229:38:@38863.4]
  assign _T_93355 = bypassInitiated_13 == 1'h0; // @[LoadQueue.scala 230:12:@38865.6]
  assign _T_93357 = prevPriorityRequest_13 == 1'h0; // @[LoadQueue.scala 230:46:@38866.6]
  assign _T_93358 = _T_93355 & _T_93357; // @[LoadQueue.scala 230:43:@38867.6]
  assign _T_93360 = dataKnown_13 == 1'h0; // @[LoadQueue.scala 230:84:@38868.6]
  assign _T_93361 = _T_93358 & _T_93360; // @[LoadQueue.scala 230:81:@38869.6]
  assign _T_93364 = storeAddrNotKnownFlagsPReg_13_0 | storeAddrNotKnownFlagsPReg_13_1; // @[LoadQueue.scala 233:86:@38872.8]
  assign _T_93365 = _T_93364 | storeAddrNotKnownFlagsPReg_13_2; // @[LoadQueue.scala 233:86:@38873.8]
  assign _T_93366 = _T_93365 | storeAddrNotKnownFlagsPReg_13_3; // @[LoadQueue.scala 233:86:@38874.8]
  assign _T_93367 = _T_93366 | storeAddrNotKnownFlagsPReg_13_4; // @[LoadQueue.scala 233:86:@38875.8]
  assign _T_93368 = _T_93367 | storeAddrNotKnownFlagsPReg_13_5; // @[LoadQueue.scala 233:86:@38876.8]
  assign _T_93369 = _T_93368 | storeAddrNotKnownFlagsPReg_13_6; // @[LoadQueue.scala 233:86:@38877.8]
  assign _T_93370 = _T_93369 | storeAddrNotKnownFlagsPReg_13_7; // @[LoadQueue.scala 233:86:@38878.8]
  assign _T_93371 = _T_93370 | storeAddrNotKnownFlagsPReg_13_8; // @[LoadQueue.scala 233:86:@38879.8]
  assign _T_93372 = _T_93371 | storeAddrNotKnownFlagsPReg_13_9; // @[LoadQueue.scala 233:86:@38880.8]
  assign _T_93373 = _T_93372 | storeAddrNotKnownFlagsPReg_13_10; // @[LoadQueue.scala 233:86:@38881.8]
  assign _T_93374 = _T_93373 | storeAddrNotKnownFlagsPReg_13_11; // @[LoadQueue.scala 233:86:@38882.8]
  assign _T_93375 = _T_93374 | storeAddrNotKnownFlagsPReg_13_12; // @[LoadQueue.scala 233:86:@38883.8]
  assign _T_93376 = _T_93375 | storeAddrNotKnownFlagsPReg_13_13; // @[LoadQueue.scala 233:86:@38884.8]
  assign _T_93377 = _T_93376 | storeAddrNotKnownFlagsPReg_13_14; // @[LoadQueue.scala 233:86:@38885.8]
  assign _T_93378 = _T_93377 | storeAddrNotKnownFlagsPReg_13_15; // @[LoadQueue.scala 233:86:@38886.8]
  assign _T_93380 = _T_93378 == 1'h0; // @[LoadQueue.scala 233:38:@38887.8]
  assign _T_93399 = _T_90074 == 1'h0; // @[LoadQueue.scala 234:11:@38904.8]
  assign _T_93400 = _T_93380 & _T_93399; // @[LoadQueue.scala 233:103:@38905.8]
  assign _GEN_2020 = _T_93361 ? _T_93400 : 1'h0; // @[LoadQueue.scala 230:110:@38870.6]
  assign loadRequest_13 = _T_93353 ? _GEN_2020 : 1'h0; // @[LoadQueue.scala 229:71:@38864.4]
  assign _T_90466 = loadRequest_13 ? 16'h2000 : _T_90465; // @[Mux.scala 31:69:@36523.4]
  assign _T_93268 = dataKnownPReg_12 == 1'h0; // @[LoadQueue.scala 229:41:@38780.4]
  assign _T_93269 = addrKnownPReg_12 & _T_93268; // @[LoadQueue.scala 229:38:@38781.4]
  assign _T_93271 = bypassInitiated_12 == 1'h0; // @[LoadQueue.scala 230:12:@38783.6]
  assign _T_93273 = prevPriorityRequest_12 == 1'h0; // @[LoadQueue.scala 230:46:@38784.6]
  assign _T_93274 = _T_93271 & _T_93273; // @[LoadQueue.scala 230:43:@38785.6]
  assign _T_93276 = dataKnown_12 == 1'h0; // @[LoadQueue.scala 230:84:@38786.6]
  assign _T_93277 = _T_93274 & _T_93276; // @[LoadQueue.scala 230:81:@38787.6]
  assign _T_93280 = storeAddrNotKnownFlagsPReg_12_0 | storeAddrNotKnownFlagsPReg_12_1; // @[LoadQueue.scala 233:86:@38790.8]
  assign _T_93281 = _T_93280 | storeAddrNotKnownFlagsPReg_12_2; // @[LoadQueue.scala 233:86:@38791.8]
  assign _T_93282 = _T_93281 | storeAddrNotKnownFlagsPReg_12_3; // @[LoadQueue.scala 233:86:@38792.8]
  assign _T_93283 = _T_93282 | storeAddrNotKnownFlagsPReg_12_4; // @[LoadQueue.scala 233:86:@38793.8]
  assign _T_93284 = _T_93283 | storeAddrNotKnownFlagsPReg_12_5; // @[LoadQueue.scala 233:86:@38794.8]
  assign _T_93285 = _T_93284 | storeAddrNotKnownFlagsPReg_12_6; // @[LoadQueue.scala 233:86:@38795.8]
  assign _T_93286 = _T_93285 | storeAddrNotKnownFlagsPReg_12_7; // @[LoadQueue.scala 233:86:@38796.8]
  assign _T_93287 = _T_93286 | storeAddrNotKnownFlagsPReg_12_8; // @[LoadQueue.scala 233:86:@38797.8]
  assign _T_93288 = _T_93287 | storeAddrNotKnownFlagsPReg_12_9; // @[LoadQueue.scala 233:86:@38798.8]
  assign _T_93289 = _T_93288 | storeAddrNotKnownFlagsPReg_12_10; // @[LoadQueue.scala 233:86:@38799.8]
  assign _T_93290 = _T_93289 | storeAddrNotKnownFlagsPReg_12_11; // @[LoadQueue.scala 233:86:@38800.8]
  assign _T_93291 = _T_93290 | storeAddrNotKnownFlagsPReg_12_12; // @[LoadQueue.scala 233:86:@38801.8]
  assign _T_93292 = _T_93291 | storeAddrNotKnownFlagsPReg_12_13; // @[LoadQueue.scala 233:86:@38802.8]
  assign _T_93293 = _T_93292 | storeAddrNotKnownFlagsPReg_12_14; // @[LoadQueue.scala 233:86:@38803.8]
  assign _T_93294 = _T_93293 | storeAddrNotKnownFlagsPReg_12_15; // @[LoadQueue.scala 233:86:@38804.8]
  assign _T_93296 = _T_93294 == 1'h0; // @[LoadQueue.scala 233:38:@38805.8]
  assign _T_93315 = _T_89938 == 1'h0; // @[LoadQueue.scala 234:11:@38822.8]
  assign _T_93316 = _T_93296 & _T_93315; // @[LoadQueue.scala 233:103:@38823.8]
  assign _GEN_2016 = _T_93277 ? _T_93316 : 1'h0; // @[LoadQueue.scala 230:110:@38788.6]
  assign loadRequest_12 = _T_93269 ? _GEN_2016 : 1'h0; // @[LoadQueue.scala 229:71:@38782.4]
  assign _T_90467 = loadRequest_12 ? 16'h1000 : _T_90466; // @[Mux.scala 31:69:@36524.4]
  assign _T_93184 = dataKnownPReg_11 == 1'h0; // @[LoadQueue.scala 229:41:@38698.4]
  assign _T_93185 = addrKnownPReg_11 & _T_93184; // @[LoadQueue.scala 229:38:@38699.4]
  assign _T_93187 = bypassInitiated_11 == 1'h0; // @[LoadQueue.scala 230:12:@38701.6]
  assign _T_93189 = prevPriorityRequest_11 == 1'h0; // @[LoadQueue.scala 230:46:@38702.6]
  assign _T_93190 = _T_93187 & _T_93189; // @[LoadQueue.scala 230:43:@38703.6]
  assign _T_93192 = dataKnown_11 == 1'h0; // @[LoadQueue.scala 230:84:@38704.6]
  assign _T_93193 = _T_93190 & _T_93192; // @[LoadQueue.scala 230:81:@38705.6]
  assign _T_93196 = storeAddrNotKnownFlagsPReg_11_0 | storeAddrNotKnownFlagsPReg_11_1; // @[LoadQueue.scala 233:86:@38708.8]
  assign _T_93197 = _T_93196 | storeAddrNotKnownFlagsPReg_11_2; // @[LoadQueue.scala 233:86:@38709.8]
  assign _T_93198 = _T_93197 | storeAddrNotKnownFlagsPReg_11_3; // @[LoadQueue.scala 233:86:@38710.8]
  assign _T_93199 = _T_93198 | storeAddrNotKnownFlagsPReg_11_4; // @[LoadQueue.scala 233:86:@38711.8]
  assign _T_93200 = _T_93199 | storeAddrNotKnownFlagsPReg_11_5; // @[LoadQueue.scala 233:86:@38712.8]
  assign _T_93201 = _T_93200 | storeAddrNotKnownFlagsPReg_11_6; // @[LoadQueue.scala 233:86:@38713.8]
  assign _T_93202 = _T_93201 | storeAddrNotKnownFlagsPReg_11_7; // @[LoadQueue.scala 233:86:@38714.8]
  assign _T_93203 = _T_93202 | storeAddrNotKnownFlagsPReg_11_8; // @[LoadQueue.scala 233:86:@38715.8]
  assign _T_93204 = _T_93203 | storeAddrNotKnownFlagsPReg_11_9; // @[LoadQueue.scala 233:86:@38716.8]
  assign _T_93205 = _T_93204 | storeAddrNotKnownFlagsPReg_11_10; // @[LoadQueue.scala 233:86:@38717.8]
  assign _T_93206 = _T_93205 | storeAddrNotKnownFlagsPReg_11_11; // @[LoadQueue.scala 233:86:@38718.8]
  assign _T_93207 = _T_93206 | storeAddrNotKnownFlagsPReg_11_12; // @[LoadQueue.scala 233:86:@38719.8]
  assign _T_93208 = _T_93207 | storeAddrNotKnownFlagsPReg_11_13; // @[LoadQueue.scala 233:86:@38720.8]
  assign _T_93209 = _T_93208 | storeAddrNotKnownFlagsPReg_11_14; // @[LoadQueue.scala 233:86:@38721.8]
  assign _T_93210 = _T_93209 | storeAddrNotKnownFlagsPReg_11_15; // @[LoadQueue.scala 233:86:@38722.8]
  assign _T_93212 = _T_93210 == 1'h0; // @[LoadQueue.scala 233:38:@38723.8]
  assign _T_93231 = _T_89802 == 1'h0; // @[LoadQueue.scala 234:11:@38740.8]
  assign _T_93232 = _T_93212 & _T_93231; // @[LoadQueue.scala 233:103:@38741.8]
  assign _GEN_2012 = _T_93193 ? _T_93232 : 1'h0; // @[LoadQueue.scala 230:110:@38706.6]
  assign loadRequest_11 = _T_93185 ? _GEN_2012 : 1'h0; // @[LoadQueue.scala 229:71:@38700.4]
  assign _T_90468 = loadRequest_11 ? 16'h800 : _T_90467; // @[Mux.scala 31:69:@36525.4]
  assign _T_93100 = dataKnownPReg_10 == 1'h0; // @[LoadQueue.scala 229:41:@38616.4]
  assign _T_93101 = addrKnownPReg_10 & _T_93100; // @[LoadQueue.scala 229:38:@38617.4]
  assign _T_93103 = bypassInitiated_10 == 1'h0; // @[LoadQueue.scala 230:12:@38619.6]
  assign _T_93105 = prevPriorityRequest_10 == 1'h0; // @[LoadQueue.scala 230:46:@38620.6]
  assign _T_93106 = _T_93103 & _T_93105; // @[LoadQueue.scala 230:43:@38621.6]
  assign _T_93108 = dataKnown_10 == 1'h0; // @[LoadQueue.scala 230:84:@38622.6]
  assign _T_93109 = _T_93106 & _T_93108; // @[LoadQueue.scala 230:81:@38623.6]
  assign _T_93112 = storeAddrNotKnownFlagsPReg_10_0 | storeAddrNotKnownFlagsPReg_10_1; // @[LoadQueue.scala 233:86:@38626.8]
  assign _T_93113 = _T_93112 | storeAddrNotKnownFlagsPReg_10_2; // @[LoadQueue.scala 233:86:@38627.8]
  assign _T_93114 = _T_93113 | storeAddrNotKnownFlagsPReg_10_3; // @[LoadQueue.scala 233:86:@38628.8]
  assign _T_93115 = _T_93114 | storeAddrNotKnownFlagsPReg_10_4; // @[LoadQueue.scala 233:86:@38629.8]
  assign _T_93116 = _T_93115 | storeAddrNotKnownFlagsPReg_10_5; // @[LoadQueue.scala 233:86:@38630.8]
  assign _T_93117 = _T_93116 | storeAddrNotKnownFlagsPReg_10_6; // @[LoadQueue.scala 233:86:@38631.8]
  assign _T_93118 = _T_93117 | storeAddrNotKnownFlagsPReg_10_7; // @[LoadQueue.scala 233:86:@38632.8]
  assign _T_93119 = _T_93118 | storeAddrNotKnownFlagsPReg_10_8; // @[LoadQueue.scala 233:86:@38633.8]
  assign _T_93120 = _T_93119 | storeAddrNotKnownFlagsPReg_10_9; // @[LoadQueue.scala 233:86:@38634.8]
  assign _T_93121 = _T_93120 | storeAddrNotKnownFlagsPReg_10_10; // @[LoadQueue.scala 233:86:@38635.8]
  assign _T_93122 = _T_93121 | storeAddrNotKnownFlagsPReg_10_11; // @[LoadQueue.scala 233:86:@38636.8]
  assign _T_93123 = _T_93122 | storeAddrNotKnownFlagsPReg_10_12; // @[LoadQueue.scala 233:86:@38637.8]
  assign _T_93124 = _T_93123 | storeAddrNotKnownFlagsPReg_10_13; // @[LoadQueue.scala 233:86:@38638.8]
  assign _T_93125 = _T_93124 | storeAddrNotKnownFlagsPReg_10_14; // @[LoadQueue.scala 233:86:@38639.8]
  assign _T_93126 = _T_93125 | storeAddrNotKnownFlagsPReg_10_15; // @[LoadQueue.scala 233:86:@38640.8]
  assign _T_93128 = _T_93126 == 1'h0; // @[LoadQueue.scala 233:38:@38641.8]
  assign _T_93147 = _T_89666 == 1'h0; // @[LoadQueue.scala 234:11:@38658.8]
  assign _T_93148 = _T_93128 & _T_93147; // @[LoadQueue.scala 233:103:@38659.8]
  assign _GEN_2008 = _T_93109 ? _T_93148 : 1'h0; // @[LoadQueue.scala 230:110:@38624.6]
  assign loadRequest_10 = _T_93101 ? _GEN_2008 : 1'h0; // @[LoadQueue.scala 229:71:@38618.4]
  assign _T_90469 = loadRequest_10 ? 16'h400 : _T_90468; // @[Mux.scala 31:69:@36526.4]
  assign _T_93016 = dataKnownPReg_9 == 1'h0; // @[LoadQueue.scala 229:41:@38534.4]
  assign _T_93017 = addrKnownPReg_9 & _T_93016; // @[LoadQueue.scala 229:38:@38535.4]
  assign _T_93019 = bypassInitiated_9 == 1'h0; // @[LoadQueue.scala 230:12:@38537.6]
  assign _T_93021 = prevPriorityRequest_9 == 1'h0; // @[LoadQueue.scala 230:46:@38538.6]
  assign _T_93022 = _T_93019 & _T_93021; // @[LoadQueue.scala 230:43:@38539.6]
  assign _T_93024 = dataKnown_9 == 1'h0; // @[LoadQueue.scala 230:84:@38540.6]
  assign _T_93025 = _T_93022 & _T_93024; // @[LoadQueue.scala 230:81:@38541.6]
  assign _T_93028 = storeAddrNotKnownFlagsPReg_9_0 | storeAddrNotKnownFlagsPReg_9_1; // @[LoadQueue.scala 233:86:@38544.8]
  assign _T_93029 = _T_93028 | storeAddrNotKnownFlagsPReg_9_2; // @[LoadQueue.scala 233:86:@38545.8]
  assign _T_93030 = _T_93029 | storeAddrNotKnownFlagsPReg_9_3; // @[LoadQueue.scala 233:86:@38546.8]
  assign _T_93031 = _T_93030 | storeAddrNotKnownFlagsPReg_9_4; // @[LoadQueue.scala 233:86:@38547.8]
  assign _T_93032 = _T_93031 | storeAddrNotKnownFlagsPReg_9_5; // @[LoadQueue.scala 233:86:@38548.8]
  assign _T_93033 = _T_93032 | storeAddrNotKnownFlagsPReg_9_6; // @[LoadQueue.scala 233:86:@38549.8]
  assign _T_93034 = _T_93033 | storeAddrNotKnownFlagsPReg_9_7; // @[LoadQueue.scala 233:86:@38550.8]
  assign _T_93035 = _T_93034 | storeAddrNotKnownFlagsPReg_9_8; // @[LoadQueue.scala 233:86:@38551.8]
  assign _T_93036 = _T_93035 | storeAddrNotKnownFlagsPReg_9_9; // @[LoadQueue.scala 233:86:@38552.8]
  assign _T_93037 = _T_93036 | storeAddrNotKnownFlagsPReg_9_10; // @[LoadQueue.scala 233:86:@38553.8]
  assign _T_93038 = _T_93037 | storeAddrNotKnownFlagsPReg_9_11; // @[LoadQueue.scala 233:86:@38554.8]
  assign _T_93039 = _T_93038 | storeAddrNotKnownFlagsPReg_9_12; // @[LoadQueue.scala 233:86:@38555.8]
  assign _T_93040 = _T_93039 | storeAddrNotKnownFlagsPReg_9_13; // @[LoadQueue.scala 233:86:@38556.8]
  assign _T_93041 = _T_93040 | storeAddrNotKnownFlagsPReg_9_14; // @[LoadQueue.scala 233:86:@38557.8]
  assign _T_93042 = _T_93041 | storeAddrNotKnownFlagsPReg_9_15; // @[LoadQueue.scala 233:86:@38558.8]
  assign _T_93044 = _T_93042 == 1'h0; // @[LoadQueue.scala 233:38:@38559.8]
  assign _T_93063 = _T_89530 == 1'h0; // @[LoadQueue.scala 234:11:@38576.8]
  assign _T_93064 = _T_93044 & _T_93063; // @[LoadQueue.scala 233:103:@38577.8]
  assign _GEN_2004 = _T_93025 ? _T_93064 : 1'h0; // @[LoadQueue.scala 230:110:@38542.6]
  assign loadRequest_9 = _T_93017 ? _GEN_2004 : 1'h0; // @[LoadQueue.scala 229:71:@38536.4]
  assign _T_90470 = loadRequest_9 ? 16'h200 : _T_90469; // @[Mux.scala 31:69:@36527.4]
  assign _T_92932 = dataKnownPReg_8 == 1'h0; // @[LoadQueue.scala 229:41:@38452.4]
  assign _T_92933 = addrKnownPReg_8 & _T_92932; // @[LoadQueue.scala 229:38:@38453.4]
  assign _T_92935 = bypassInitiated_8 == 1'h0; // @[LoadQueue.scala 230:12:@38455.6]
  assign _T_92937 = prevPriorityRequest_8 == 1'h0; // @[LoadQueue.scala 230:46:@38456.6]
  assign _T_92938 = _T_92935 & _T_92937; // @[LoadQueue.scala 230:43:@38457.6]
  assign _T_92940 = dataKnown_8 == 1'h0; // @[LoadQueue.scala 230:84:@38458.6]
  assign _T_92941 = _T_92938 & _T_92940; // @[LoadQueue.scala 230:81:@38459.6]
  assign _T_92944 = storeAddrNotKnownFlagsPReg_8_0 | storeAddrNotKnownFlagsPReg_8_1; // @[LoadQueue.scala 233:86:@38462.8]
  assign _T_92945 = _T_92944 | storeAddrNotKnownFlagsPReg_8_2; // @[LoadQueue.scala 233:86:@38463.8]
  assign _T_92946 = _T_92945 | storeAddrNotKnownFlagsPReg_8_3; // @[LoadQueue.scala 233:86:@38464.8]
  assign _T_92947 = _T_92946 | storeAddrNotKnownFlagsPReg_8_4; // @[LoadQueue.scala 233:86:@38465.8]
  assign _T_92948 = _T_92947 | storeAddrNotKnownFlagsPReg_8_5; // @[LoadQueue.scala 233:86:@38466.8]
  assign _T_92949 = _T_92948 | storeAddrNotKnownFlagsPReg_8_6; // @[LoadQueue.scala 233:86:@38467.8]
  assign _T_92950 = _T_92949 | storeAddrNotKnownFlagsPReg_8_7; // @[LoadQueue.scala 233:86:@38468.8]
  assign _T_92951 = _T_92950 | storeAddrNotKnownFlagsPReg_8_8; // @[LoadQueue.scala 233:86:@38469.8]
  assign _T_92952 = _T_92951 | storeAddrNotKnownFlagsPReg_8_9; // @[LoadQueue.scala 233:86:@38470.8]
  assign _T_92953 = _T_92952 | storeAddrNotKnownFlagsPReg_8_10; // @[LoadQueue.scala 233:86:@38471.8]
  assign _T_92954 = _T_92953 | storeAddrNotKnownFlagsPReg_8_11; // @[LoadQueue.scala 233:86:@38472.8]
  assign _T_92955 = _T_92954 | storeAddrNotKnownFlagsPReg_8_12; // @[LoadQueue.scala 233:86:@38473.8]
  assign _T_92956 = _T_92955 | storeAddrNotKnownFlagsPReg_8_13; // @[LoadQueue.scala 233:86:@38474.8]
  assign _T_92957 = _T_92956 | storeAddrNotKnownFlagsPReg_8_14; // @[LoadQueue.scala 233:86:@38475.8]
  assign _T_92958 = _T_92957 | storeAddrNotKnownFlagsPReg_8_15; // @[LoadQueue.scala 233:86:@38476.8]
  assign _T_92960 = _T_92958 == 1'h0; // @[LoadQueue.scala 233:38:@38477.8]
  assign _T_92979 = _T_89394 == 1'h0; // @[LoadQueue.scala 234:11:@38494.8]
  assign _T_92980 = _T_92960 & _T_92979; // @[LoadQueue.scala 233:103:@38495.8]
  assign _GEN_2000 = _T_92941 ? _T_92980 : 1'h0; // @[LoadQueue.scala 230:110:@38460.6]
  assign loadRequest_8 = _T_92933 ? _GEN_2000 : 1'h0; // @[LoadQueue.scala 229:71:@38454.4]
  assign _T_90471 = loadRequest_8 ? 16'h100 : _T_90470; // @[Mux.scala 31:69:@36528.4]
  assign _T_92848 = dataKnownPReg_7 == 1'h0; // @[LoadQueue.scala 229:41:@38370.4]
  assign _T_92849 = addrKnownPReg_7 & _T_92848; // @[LoadQueue.scala 229:38:@38371.4]
  assign _T_92851 = bypassInitiated_7 == 1'h0; // @[LoadQueue.scala 230:12:@38373.6]
  assign _T_92853 = prevPriorityRequest_7 == 1'h0; // @[LoadQueue.scala 230:46:@38374.6]
  assign _T_92854 = _T_92851 & _T_92853; // @[LoadQueue.scala 230:43:@38375.6]
  assign _T_92856 = dataKnown_7 == 1'h0; // @[LoadQueue.scala 230:84:@38376.6]
  assign _T_92857 = _T_92854 & _T_92856; // @[LoadQueue.scala 230:81:@38377.6]
  assign _T_92860 = storeAddrNotKnownFlagsPReg_7_0 | storeAddrNotKnownFlagsPReg_7_1; // @[LoadQueue.scala 233:86:@38380.8]
  assign _T_92861 = _T_92860 | storeAddrNotKnownFlagsPReg_7_2; // @[LoadQueue.scala 233:86:@38381.8]
  assign _T_92862 = _T_92861 | storeAddrNotKnownFlagsPReg_7_3; // @[LoadQueue.scala 233:86:@38382.8]
  assign _T_92863 = _T_92862 | storeAddrNotKnownFlagsPReg_7_4; // @[LoadQueue.scala 233:86:@38383.8]
  assign _T_92864 = _T_92863 | storeAddrNotKnownFlagsPReg_7_5; // @[LoadQueue.scala 233:86:@38384.8]
  assign _T_92865 = _T_92864 | storeAddrNotKnownFlagsPReg_7_6; // @[LoadQueue.scala 233:86:@38385.8]
  assign _T_92866 = _T_92865 | storeAddrNotKnownFlagsPReg_7_7; // @[LoadQueue.scala 233:86:@38386.8]
  assign _T_92867 = _T_92866 | storeAddrNotKnownFlagsPReg_7_8; // @[LoadQueue.scala 233:86:@38387.8]
  assign _T_92868 = _T_92867 | storeAddrNotKnownFlagsPReg_7_9; // @[LoadQueue.scala 233:86:@38388.8]
  assign _T_92869 = _T_92868 | storeAddrNotKnownFlagsPReg_7_10; // @[LoadQueue.scala 233:86:@38389.8]
  assign _T_92870 = _T_92869 | storeAddrNotKnownFlagsPReg_7_11; // @[LoadQueue.scala 233:86:@38390.8]
  assign _T_92871 = _T_92870 | storeAddrNotKnownFlagsPReg_7_12; // @[LoadQueue.scala 233:86:@38391.8]
  assign _T_92872 = _T_92871 | storeAddrNotKnownFlagsPReg_7_13; // @[LoadQueue.scala 233:86:@38392.8]
  assign _T_92873 = _T_92872 | storeAddrNotKnownFlagsPReg_7_14; // @[LoadQueue.scala 233:86:@38393.8]
  assign _T_92874 = _T_92873 | storeAddrNotKnownFlagsPReg_7_15; // @[LoadQueue.scala 233:86:@38394.8]
  assign _T_92876 = _T_92874 == 1'h0; // @[LoadQueue.scala 233:38:@38395.8]
  assign _T_92895 = _T_89258 == 1'h0; // @[LoadQueue.scala 234:11:@38412.8]
  assign _T_92896 = _T_92876 & _T_92895; // @[LoadQueue.scala 233:103:@38413.8]
  assign _GEN_1996 = _T_92857 ? _T_92896 : 1'h0; // @[LoadQueue.scala 230:110:@38378.6]
  assign loadRequest_7 = _T_92849 ? _GEN_1996 : 1'h0; // @[LoadQueue.scala 229:71:@38372.4]
  assign _T_90472 = loadRequest_7 ? 16'h80 : _T_90471; // @[Mux.scala 31:69:@36529.4]
  assign _T_92764 = dataKnownPReg_6 == 1'h0; // @[LoadQueue.scala 229:41:@38288.4]
  assign _T_92765 = addrKnownPReg_6 & _T_92764; // @[LoadQueue.scala 229:38:@38289.4]
  assign _T_92767 = bypassInitiated_6 == 1'h0; // @[LoadQueue.scala 230:12:@38291.6]
  assign _T_92769 = prevPriorityRequest_6 == 1'h0; // @[LoadQueue.scala 230:46:@38292.6]
  assign _T_92770 = _T_92767 & _T_92769; // @[LoadQueue.scala 230:43:@38293.6]
  assign _T_92772 = dataKnown_6 == 1'h0; // @[LoadQueue.scala 230:84:@38294.6]
  assign _T_92773 = _T_92770 & _T_92772; // @[LoadQueue.scala 230:81:@38295.6]
  assign _T_92776 = storeAddrNotKnownFlagsPReg_6_0 | storeAddrNotKnownFlagsPReg_6_1; // @[LoadQueue.scala 233:86:@38298.8]
  assign _T_92777 = _T_92776 | storeAddrNotKnownFlagsPReg_6_2; // @[LoadQueue.scala 233:86:@38299.8]
  assign _T_92778 = _T_92777 | storeAddrNotKnownFlagsPReg_6_3; // @[LoadQueue.scala 233:86:@38300.8]
  assign _T_92779 = _T_92778 | storeAddrNotKnownFlagsPReg_6_4; // @[LoadQueue.scala 233:86:@38301.8]
  assign _T_92780 = _T_92779 | storeAddrNotKnownFlagsPReg_6_5; // @[LoadQueue.scala 233:86:@38302.8]
  assign _T_92781 = _T_92780 | storeAddrNotKnownFlagsPReg_6_6; // @[LoadQueue.scala 233:86:@38303.8]
  assign _T_92782 = _T_92781 | storeAddrNotKnownFlagsPReg_6_7; // @[LoadQueue.scala 233:86:@38304.8]
  assign _T_92783 = _T_92782 | storeAddrNotKnownFlagsPReg_6_8; // @[LoadQueue.scala 233:86:@38305.8]
  assign _T_92784 = _T_92783 | storeAddrNotKnownFlagsPReg_6_9; // @[LoadQueue.scala 233:86:@38306.8]
  assign _T_92785 = _T_92784 | storeAddrNotKnownFlagsPReg_6_10; // @[LoadQueue.scala 233:86:@38307.8]
  assign _T_92786 = _T_92785 | storeAddrNotKnownFlagsPReg_6_11; // @[LoadQueue.scala 233:86:@38308.8]
  assign _T_92787 = _T_92786 | storeAddrNotKnownFlagsPReg_6_12; // @[LoadQueue.scala 233:86:@38309.8]
  assign _T_92788 = _T_92787 | storeAddrNotKnownFlagsPReg_6_13; // @[LoadQueue.scala 233:86:@38310.8]
  assign _T_92789 = _T_92788 | storeAddrNotKnownFlagsPReg_6_14; // @[LoadQueue.scala 233:86:@38311.8]
  assign _T_92790 = _T_92789 | storeAddrNotKnownFlagsPReg_6_15; // @[LoadQueue.scala 233:86:@38312.8]
  assign _T_92792 = _T_92790 == 1'h0; // @[LoadQueue.scala 233:38:@38313.8]
  assign _T_92811 = _T_89122 == 1'h0; // @[LoadQueue.scala 234:11:@38330.8]
  assign _T_92812 = _T_92792 & _T_92811; // @[LoadQueue.scala 233:103:@38331.8]
  assign _GEN_1992 = _T_92773 ? _T_92812 : 1'h0; // @[LoadQueue.scala 230:110:@38296.6]
  assign loadRequest_6 = _T_92765 ? _GEN_1992 : 1'h0; // @[LoadQueue.scala 229:71:@38290.4]
  assign _T_90473 = loadRequest_6 ? 16'h40 : _T_90472; // @[Mux.scala 31:69:@36530.4]
  assign _T_92680 = dataKnownPReg_5 == 1'h0; // @[LoadQueue.scala 229:41:@38206.4]
  assign _T_92681 = addrKnownPReg_5 & _T_92680; // @[LoadQueue.scala 229:38:@38207.4]
  assign _T_92683 = bypassInitiated_5 == 1'h0; // @[LoadQueue.scala 230:12:@38209.6]
  assign _T_92685 = prevPriorityRequest_5 == 1'h0; // @[LoadQueue.scala 230:46:@38210.6]
  assign _T_92686 = _T_92683 & _T_92685; // @[LoadQueue.scala 230:43:@38211.6]
  assign _T_92688 = dataKnown_5 == 1'h0; // @[LoadQueue.scala 230:84:@38212.6]
  assign _T_92689 = _T_92686 & _T_92688; // @[LoadQueue.scala 230:81:@38213.6]
  assign _T_92692 = storeAddrNotKnownFlagsPReg_5_0 | storeAddrNotKnownFlagsPReg_5_1; // @[LoadQueue.scala 233:86:@38216.8]
  assign _T_92693 = _T_92692 | storeAddrNotKnownFlagsPReg_5_2; // @[LoadQueue.scala 233:86:@38217.8]
  assign _T_92694 = _T_92693 | storeAddrNotKnownFlagsPReg_5_3; // @[LoadQueue.scala 233:86:@38218.8]
  assign _T_92695 = _T_92694 | storeAddrNotKnownFlagsPReg_5_4; // @[LoadQueue.scala 233:86:@38219.8]
  assign _T_92696 = _T_92695 | storeAddrNotKnownFlagsPReg_5_5; // @[LoadQueue.scala 233:86:@38220.8]
  assign _T_92697 = _T_92696 | storeAddrNotKnownFlagsPReg_5_6; // @[LoadQueue.scala 233:86:@38221.8]
  assign _T_92698 = _T_92697 | storeAddrNotKnownFlagsPReg_5_7; // @[LoadQueue.scala 233:86:@38222.8]
  assign _T_92699 = _T_92698 | storeAddrNotKnownFlagsPReg_5_8; // @[LoadQueue.scala 233:86:@38223.8]
  assign _T_92700 = _T_92699 | storeAddrNotKnownFlagsPReg_5_9; // @[LoadQueue.scala 233:86:@38224.8]
  assign _T_92701 = _T_92700 | storeAddrNotKnownFlagsPReg_5_10; // @[LoadQueue.scala 233:86:@38225.8]
  assign _T_92702 = _T_92701 | storeAddrNotKnownFlagsPReg_5_11; // @[LoadQueue.scala 233:86:@38226.8]
  assign _T_92703 = _T_92702 | storeAddrNotKnownFlagsPReg_5_12; // @[LoadQueue.scala 233:86:@38227.8]
  assign _T_92704 = _T_92703 | storeAddrNotKnownFlagsPReg_5_13; // @[LoadQueue.scala 233:86:@38228.8]
  assign _T_92705 = _T_92704 | storeAddrNotKnownFlagsPReg_5_14; // @[LoadQueue.scala 233:86:@38229.8]
  assign _T_92706 = _T_92705 | storeAddrNotKnownFlagsPReg_5_15; // @[LoadQueue.scala 233:86:@38230.8]
  assign _T_92708 = _T_92706 == 1'h0; // @[LoadQueue.scala 233:38:@38231.8]
  assign _T_92727 = _T_88986 == 1'h0; // @[LoadQueue.scala 234:11:@38248.8]
  assign _T_92728 = _T_92708 & _T_92727; // @[LoadQueue.scala 233:103:@38249.8]
  assign _GEN_1988 = _T_92689 ? _T_92728 : 1'h0; // @[LoadQueue.scala 230:110:@38214.6]
  assign loadRequest_5 = _T_92681 ? _GEN_1988 : 1'h0; // @[LoadQueue.scala 229:71:@38208.4]
  assign _T_90474 = loadRequest_5 ? 16'h20 : _T_90473; // @[Mux.scala 31:69:@36531.4]
  assign _T_92596 = dataKnownPReg_4 == 1'h0; // @[LoadQueue.scala 229:41:@38124.4]
  assign _T_92597 = addrKnownPReg_4 & _T_92596; // @[LoadQueue.scala 229:38:@38125.4]
  assign _T_92599 = bypassInitiated_4 == 1'h0; // @[LoadQueue.scala 230:12:@38127.6]
  assign _T_92601 = prevPriorityRequest_4 == 1'h0; // @[LoadQueue.scala 230:46:@38128.6]
  assign _T_92602 = _T_92599 & _T_92601; // @[LoadQueue.scala 230:43:@38129.6]
  assign _T_92604 = dataKnown_4 == 1'h0; // @[LoadQueue.scala 230:84:@38130.6]
  assign _T_92605 = _T_92602 & _T_92604; // @[LoadQueue.scala 230:81:@38131.6]
  assign _T_92608 = storeAddrNotKnownFlagsPReg_4_0 | storeAddrNotKnownFlagsPReg_4_1; // @[LoadQueue.scala 233:86:@38134.8]
  assign _T_92609 = _T_92608 | storeAddrNotKnownFlagsPReg_4_2; // @[LoadQueue.scala 233:86:@38135.8]
  assign _T_92610 = _T_92609 | storeAddrNotKnownFlagsPReg_4_3; // @[LoadQueue.scala 233:86:@38136.8]
  assign _T_92611 = _T_92610 | storeAddrNotKnownFlagsPReg_4_4; // @[LoadQueue.scala 233:86:@38137.8]
  assign _T_92612 = _T_92611 | storeAddrNotKnownFlagsPReg_4_5; // @[LoadQueue.scala 233:86:@38138.8]
  assign _T_92613 = _T_92612 | storeAddrNotKnownFlagsPReg_4_6; // @[LoadQueue.scala 233:86:@38139.8]
  assign _T_92614 = _T_92613 | storeAddrNotKnownFlagsPReg_4_7; // @[LoadQueue.scala 233:86:@38140.8]
  assign _T_92615 = _T_92614 | storeAddrNotKnownFlagsPReg_4_8; // @[LoadQueue.scala 233:86:@38141.8]
  assign _T_92616 = _T_92615 | storeAddrNotKnownFlagsPReg_4_9; // @[LoadQueue.scala 233:86:@38142.8]
  assign _T_92617 = _T_92616 | storeAddrNotKnownFlagsPReg_4_10; // @[LoadQueue.scala 233:86:@38143.8]
  assign _T_92618 = _T_92617 | storeAddrNotKnownFlagsPReg_4_11; // @[LoadQueue.scala 233:86:@38144.8]
  assign _T_92619 = _T_92618 | storeAddrNotKnownFlagsPReg_4_12; // @[LoadQueue.scala 233:86:@38145.8]
  assign _T_92620 = _T_92619 | storeAddrNotKnownFlagsPReg_4_13; // @[LoadQueue.scala 233:86:@38146.8]
  assign _T_92621 = _T_92620 | storeAddrNotKnownFlagsPReg_4_14; // @[LoadQueue.scala 233:86:@38147.8]
  assign _T_92622 = _T_92621 | storeAddrNotKnownFlagsPReg_4_15; // @[LoadQueue.scala 233:86:@38148.8]
  assign _T_92624 = _T_92622 == 1'h0; // @[LoadQueue.scala 233:38:@38149.8]
  assign _T_92643 = _T_88850 == 1'h0; // @[LoadQueue.scala 234:11:@38166.8]
  assign _T_92644 = _T_92624 & _T_92643; // @[LoadQueue.scala 233:103:@38167.8]
  assign _GEN_1984 = _T_92605 ? _T_92644 : 1'h0; // @[LoadQueue.scala 230:110:@38132.6]
  assign loadRequest_4 = _T_92597 ? _GEN_1984 : 1'h0; // @[LoadQueue.scala 229:71:@38126.4]
  assign _T_90475 = loadRequest_4 ? 16'h10 : _T_90474; // @[Mux.scala 31:69:@36532.4]
  assign _T_92512 = dataKnownPReg_3 == 1'h0; // @[LoadQueue.scala 229:41:@38042.4]
  assign _T_92513 = addrKnownPReg_3 & _T_92512; // @[LoadQueue.scala 229:38:@38043.4]
  assign _T_92515 = bypassInitiated_3 == 1'h0; // @[LoadQueue.scala 230:12:@38045.6]
  assign _T_92517 = prevPriorityRequest_3 == 1'h0; // @[LoadQueue.scala 230:46:@38046.6]
  assign _T_92518 = _T_92515 & _T_92517; // @[LoadQueue.scala 230:43:@38047.6]
  assign _T_92520 = dataKnown_3 == 1'h0; // @[LoadQueue.scala 230:84:@38048.6]
  assign _T_92521 = _T_92518 & _T_92520; // @[LoadQueue.scala 230:81:@38049.6]
  assign _T_92524 = storeAddrNotKnownFlagsPReg_3_0 | storeAddrNotKnownFlagsPReg_3_1; // @[LoadQueue.scala 233:86:@38052.8]
  assign _T_92525 = _T_92524 | storeAddrNotKnownFlagsPReg_3_2; // @[LoadQueue.scala 233:86:@38053.8]
  assign _T_92526 = _T_92525 | storeAddrNotKnownFlagsPReg_3_3; // @[LoadQueue.scala 233:86:@38054.8]
  assign _T_92527 = _T_92526 | storeAddrNotKnownFlagsPReg_3_4; // @[LoadQueue.scala 233:86:@38055.8]
  assign _T_92528 = _T_92527 | storeAddrNotKnownFlagsPReg_3_5; // @[LoadQueue.scala 233:86:@38056.8]
  assign _T_92529 = _T_92528 | storeAddrNotKnownFlagsPReg_3_6; // @[LoadQueue.scala 233:86:@38057.8]
  assign _T_92530 = _T_92529 | storeAddrNotKnownFlagsPReg_3_7; // @[LoadQueue.scala 233:86:@38058.8]
  assign _T_92531 = _T_92530 | storeAddrNotKnownFlagsPReg_3_8; // @[LoadQueue.scala 233:86:@38059.8]
  assign _T_92532 = _T_92531 | storeAddrNotKnownFlagsPReg_3_9; // @[LoadQueue.scala 233:86:@38060.8]
  assign _T_92533 = _T_92532 | storeAddrNotKnownFlagsPReg_3_10; // @[LoadQueue.scala 233:86:@38061.8]
  assign _T_92534 = _T_92533 | storeAddrNotKnownFlagsPReg_3_11; // @[LoadQueue.scala 233:86:@38062.8]
  assign _T_92535 = _T_92534 | storeAddrNotKnownFlagsPReg_3_12; // @[LoadQueue.scala 233:86:@38063.8]
  assign _T_92536 = _T_92535 | storeAddrNotKnownFlagsPReg_3_13; // @[LoadQueue.scala 233:86:@38064.8]
  assign _T_92537 = _T_92536 | storeAddrNotKnownFlagsPReg_3_14; // @[LoadQueue.scala 233:86:@38065.8]
  assign _T_92538 = _T_92537 | storeAddrNotKnownFlagsPReg_3_15; // @[LoadQueue.scala 233:86:@38066.8]
  assign _T_92540 = _T_92538 == 1'h0; // @[LoadQueue.scala 233:38:@38067.8]
  assign _T_92559 = _T_88714 == 1'h0; // @[LoadQueue.scala 234:11:@38084.8]
  assign _T_92560 = _T_92540 & _T_92559; // @[LoadQueue.scala 233:103:@38085.8]
  assign _GEN_1980 = _T_92521 ? _T_92560 : 1'h0; // @[LoadQueue.scala 230:110:@38050.6]
  assign loadRequest_3 = _T_92513 ? _GEN_1980 : 1'h0; // @[LoadQueue.scala 229:71:@38044.4]
  assign _T_90476 = loadRequest_3 ? 16'h8 : _T_90475; // @[Mux.scala 31:69:@36533.4]
  assign _T_92428 = dataKnownPReg_2 == 1'h0; // @[LoadQueue.scala 229:41:@37960.4]
  assign _T_92429 = addrKnownPReg_2 & _T_92428; // @[LoadQueue.scala 229:38:@37961.4]
  assign _T_92431 = bypassInitiated_2 == 1'h0; // @[LoadQueue.scala 230:12:@37963.6]
  assign _T_92433 = prevPriorityRequest_2 == 1'h0; // @[LoadQueue.scala 230:46:@37964.6]
  assign _T_92434 = _T_92431 & _T_92433; // @[LoadQueue.scala 230:43:@37965.6]
  assign _T_92436 = dataKnown_2 == 1'h0; // @[LoadQueue.scala 230:84:@37966.6]
  assign _T_92437 = _T_92434 & _T_92436; // @[LoadQueue.scala 230:81:@37967.6]
  assign _T_92440 = storeAddrNotKnownFlagsPReg_2_0 | storeAddrNotKnownFlagsPReg_2_1; // @[LoadQueue.scala 233:86:@37970.8]
  assign _T_92441 = _T_92440 | storeAddrNotKnownFlagsPReg_2_2; // @[LoadQueue.scala 233:86:@37971.8]
  assign _T_92442 = _T_92441 | storeAddrNotKnownFlagsPReg_2_3; // @[LoadQueue.scala 233:86:@37972.8]
  assign _T_92443 = _T_92442 | storeAddrNotKnownFlagsPReg_2_4; // @[LoadQueue.scala 233:86:@37973.8]
  assign _T_92444 = _T_92443 | storeAddrNotKnownFlagsPReg_2_5; // @[LoadQueue.scala 233:86:@37974.8]
  assign _T_92445 = _T_92444 | storeAddrNotKnownFlagsPReg_2_6; // @[LoadQueue.scala 233:86:@37975.8]
  assign _T_92446 = _T_92445 | storeAddrNotKnownFlagsPReg_2_7; // @[LoadQueue.scala 233:86:@37976.8]
  assign _T_92447 = _T_92446 | storeAddrNotKnownFlagsPReg_2_8; // @[LoadQueue.scala 233:86:@37977.8]
  assign _T_92448 = _T_92447 | storeAddrNotKnownFlagsPReg_2_9; // @[LoadQueue.scala 233:86:@37978.8]
  assign _T_92449 = _T_92448 | storeAddrNotKnownFlagsPReg_2_10; // @[LoadQueue.scala 233:86:@37979.8]
  assign _T_92450 = _T_92449 | storeAddrNotKnownFlagsPReg_2_11; // @[LoadQueue.scala 233:86:@37980.8]
  assign _T_92451 = _T_92450 | storeAddrNotKnownFlagsPReg_2_12; // @[LoadQueue.scala 233:86:@37981.8]
  assign _T_92452 = _T_92451 | storeAddrNotKnownFlagsPReg_2_13; // @[LoadQueue.scala 233:86:@37982.8]
  assign _T_92453 = _T_92452 | storeAddrNotKnownFlagsPReg_2_14; // @[LoadQueue.scala 233:86:@37983.8]
  assign _T_92454 = _T_92453 | storeAddrNotKnownFlagsPReg_2_15; // @[LoadQueue.scala 233:86:@37984.8]
  assign _T_92456 = _T_92454 == 1'h0; // @[LoadQueue.scala 233:38:@37985.8]
  assign _T_92475 = _T_88578 == 1'h0; // @[LoadQueue.scala 234:11:@38002.8]
  assign _T_92476 = _T_92456 & _T_92475; // @[LoadQueue.scala 233:103:@38003.8]
  assign _GEN_1976 = _T_92437 ? _T_92476 : 1'h0; // @[LoadQueue.scala 230:110:@37968.6]
  assign loadRequest_2 = _T_92429 ? _GEN_1976 : 1'h0; // @[LoadQueue.scala 229:71:@37962.4]
  assign _T_90477 = loadRequest_2 ? 16'h4 : _T_90476; // @[Mux.scala 31:69:@36534.4]
  assign _T_92344 = dataKnownPReg_1 == 1'h0; // @[LoadQueue.scala 229:41:@37878.4]
  assign _T_92345 = addrKnownPReg_1 & _T_92344; // @[LoadQueue.scala 229:38:@37879.4]
  assign _T_92347 = bypassInitiated_1 == 1'h0; // @[LoadQueue.scala 230:12:@37881.6]
  assign _T_92349 = prevPriorityRequest_1 == 1'h0; // @[LoadQueue.scala 230:46:@37882.6]
  assign _T_92350 = _T_92347 & _T_92349; // @[LoadQueue.scala 230:43:@37883.6]
  assign _T_92352 = dataKnown_1 == 1'h0; // @[LoadQueue.scala 230:84:@37884.6]
  assign _T_92353 = _T_92350 & _T_92352; // @[LoadQueue.scala 230:81:@37885.6]
  assign _T_92356 = storeAddrNotKnownFlagsPReg_1_0 | storeAddrNotKnownFlagsPReg_1_1; // @[LoadQueue.scala 233:86:@37888.8]
  assign _T_92357 = _T_92356 | storeAddrNotKnownFlagsPReg_1_2; // @[LoadQueue.scala 233:86:@37889.8]
  assign _T_92358 = _T_92357 | storeAddrNotKnownFlagsPReg_1_3; // @[LoadQueue.scala 233:86:@37890.8]
  assign _T_92359 = _T_92358 | storeAddrNotKnownFlagsPReg_1_4; // @[LoadQueue.scala 233:86:@37891.8]
  assign _T_92360 = _T_92359 | storeAddrNotKnownFlagsPReg_1_5; // @[LoadQueue.scala 233:86:@37892.8]
  assign _T_92361 = _T_92360 | storeAddrNotKnownFlagsPReg_1_6; // @[LoadQueue.scala 233:86:@37893.8]
  assign _T_92362 = _T_92361 | storeAddrNotKnownFlagsPReg_1_7; // @[LoadQueue.scala 233:86:@37894.8]
  assign _T_92363 = _T_92362 | storeAddrNotKnownFlagsPReg_1_8; // @[LoadQueue.scala 233:86:@37895.8]
  assign _T_92364 = _T_92363 | storeAddrNotKnownFlagsPReg_1_9; // @[LoadQueue.scala 233:86:@37896.8]
  assign _T_92365 = _T_92364 | storeAddrNotKnownFlagsPReg_1_10; // @[LoadQueue.scala 233:86:@37897.8]
  assign _T_92366 = _T_92365 | storeAddrNotKnownFlagsPReg_1_11; // @[LoadQueue.scala 233:86:@37898.8]
  assign _T_92367 = _T_92366 | storeAddrNotKnownFlagsPReg_1_12; // @[LoadQueue.scala 233:86:@37899.8]
  assign _T_92368 = _T_92367 | storeAddrNotKnownFlagsPReg_1_13; // @[LoadQueue.scala 233:86:@37900.8]
  assign _T_92369 = _T_92368 | storeAddrNotKnownFlagsPReg_1_14; // @[LoadQueue.scala 233:86:@37901.8]
  assign _T_92370 = _T_92369 | storeAddrNotKnownFlagsPReg_1_15; // @[LoadQueue.scala 233:86:@37902.8]
  assign _T_92372 = _T_92370 == 1'h0; // @[LoadQueue.scala 233:38:@37903.8]
  assign _T_92391 = _T_88442 == 1'h0; // @[LoadQueue.scala 234:11:@37920.8]
  assign _T_92392 = _T_92372 & _T_92391; // @[LoadQueue.scala 233:103:@37921.8]
  assign _GEN_1972 = _T_92353 ? _T_92392 : 1'h0; // @[LoadQueue.scala 230:110:@37886.6]
  assign loadRequest_1 = _T_92345 ? _GEN_1972 : 1'h0; // @[LoadQueue.scala 229:71:@37880.4]
  assign _T_90478 = loadRequest_1 ? 16'h2 : _T_90477; // @[Mux.scala 31:69:@36535.4]
  assign _T_92260 = dataKnownPReg_0 == 1'h0; // @[LoadQueue.scala 229:41:@37796.4]
  assign _T_92261 = addrKnownPReg_0 & _T_92260; // @[LoadQueue.scala 229:38:@37797.4]
  assign _T_92263 = bypassInitiated_0 == 1'h0; // @[LoadQueue.scala 230:12:@37799.6]
  assign _T_92265 = prevPriorityRequest_0 == 1'h0; // @[LoadQueue.scala 230:46:@37800.6]
  assign _T_92266 = _T_92263 & _T_92265; // @[LoadQueue.scala 230:43:@37801.6]
  assign _T_92268 = dataKnown_0 == 1'h0; // @[LoadQueue.scala 230:84:@37802.6]
  assign _T_92269 = _T_92266 & _T_92268; // @[LoadQueue.scala 230:81:@37803.6]
  assign _T_92272 = storeAddrNotKnownFlagsPReg_0_0 | storeAddrNotKnownFlagsPReg_0_1; // @[LoadQueue.scala 233:86:@37806.8]
  assign _T_92273 = _T_92272 | storeAddrNotKnownFlagsPReg_0_2; // @[LoadQueue.scala 233:86:@37807.8]
  assign _T_92274 = _T_92273 | storeAddrNotKnownFlagsPReg_0_3; // @[LoadQueue.scala 233:86:@37808.8]
  assign _T_92275 = _T_92274 | storeAddrNotKnownFlagsPReg_0_4; // @[LoadQueue.scala 233:86:@37809.8]
  assign _T_92276 = _T_92275 | storeAddrNotKnownFlagsPReg_0_5; // @[LoadQueue.scala 233:86:@37810.8]
  assign _T_92277 = _T_92276 | storeAddrNotKnownFlagsPReg_0_6; // @[LoadQueue.scala 233:86:@37811.8]
  assign _T_92278 = _T_92277 | storeAddrNotKnownFlagsPReg_0_7; // @[LoadQueue.scala 233:86:@37812.8]
  assign _T_92279 = _T_92278 | storeAddrNotKnownFlagsPReg_0_8; // @[LoadQueue.scala 233:86:@37813.8]
  assign _T_92280 = _T_92279 | storeAddrNotKnownFlagsPReg_0_9; // @[LoadQueue.scala 233:86:@37814.8]
  assign _T_92281 = _T_92280 | storeAddrNotKnownFlagsPReg_0_10; // @[LoadQueue.scala 233:86:@37815.8]
  assign _T_92282 = _T_92281 | storeAddrNotKnownFlagsPReg_0_11; // @[LoadQueue.scala 233:86:@37816.8]
  assign _T_92283 = _T_92282 | storeAddrNotKnownFlagsPReg_0_12; // @[LoadQueue.scala 233:86:@37817.8]
  assign _T_92284 = _T_92283 | storeAddrNotKnownFlagsPReg_0_13; // @[LoadQueue.scala 233:86:@37818.8]
  assign _T_92285 = _T_92284 | storeAddrNotKnownFlagsPReg_0_14; // @[LoadQueue.scala 233:86:@37819.8]
  assign _T_92286 = _T_92285 | storeAddrNotKnownFlagsPReg_0_15; // @[LoadQueue.scala 233:86:@37820.8]
  assign _T_92288 = _T_92286 == 1'h0; // @[LoadQueue.scala 233:38:@37821.8]
  assign _T_92307 = _T_88306 == 1'h0; // @[LoadQueue.scala 234:11:@37838.8]
  assign _T_92308 = _T_92288 & _T_92307; // @[LoadQueue.scala 233:103:@37839.8]
  assign _GEN_1968 = _T_92269 ? _T_92308 : 1'h0; // @[LoadQueue.scala 230:110:@37804.6]
  assign loadRequest_0 = _T_92261 ? _GEN_1968 : 1'h0; // @[LoadQueue.scala 229:71:@37798.4]
  assign _T_90479 = loadRequest_0 ? 16'h1 : _T_90478; // @[Mux.scala 31:69:@36536.4]
  assign _T_90480 = _T_90479[0]; // @[OneHot.scala 66:30:@36537.4]
  assign _T_90481 = _T_90479[1]; // @[OneHot.scala 66:30:@36538.4]
  assign _T_90482 = _T_90479[2]; // @[OneHot.scala 66:30:@36539.4]
  assign _T_90483 = _T_90479[3]; // @[OneHot.scala 66:30:@36540.4]
  assign _T_90484 = _T_90479[4]; // @[OneHot.scala 66:30:@36541.4]
  assign _T_90485 = _T_90479[5]; // @[OneHot.scala 66:30:@36542.4]
  assign _T_90486 = _T_90479[6]; // @[OneHot.scala 66:30:@36543.4]
  assign _T_90487 = _T_90479[7]; // @[OneHot.scala 66:30:@36544.4]
  assign _T_90488 = _T_90479[8]; // @[OneHot.scala 66:30:@36545.4]
  assign _T_90489 = _T_90479[9]; // @[OneHot.scala 66:30:@36546.4]
  assign _T_90490 = _T_90479[10]; // @[OneHot.scala 66:30:@36547.4]
  assign _T_90491 = _T_90479[11]; // @[OneHot.scala 66:30:@36548.4]
  assign _T_90492 = _T_90479[12]; // @[OneHot.scala 66:30:@36549.4]
  assign _T_90493 = _T_90479[13]; // @[OneHot.scala 66:30:@36550.4]
  assign _T_90494 = _T_90479[14]; // @[OneHot.scala 66:30:@36551.4]
  assign _T_90495 = _T_90479[15]; // @[OneHot.scala 66:30:@36552.4]
  assign _T_90536 = loadRequest_0 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36570.4]
  assign _T_90537 = loadRequest_15 ? 16'h4000 : _T_90536; // @[Mux.scala 31:69:@36571.4]
  assign _T_90538 = loadRequest_14 ? 16'h2000 : _T_90537; // @[Mux.scala 31:69:@36572.4]
  assign _T_90539 = loadRequest_13 ? 16'h1000 : _T_90538; // @[Mux.scala 31:69:@36573.4]
  assign _T_90540 = loadRequest_12 ? 16'h800 : _T_90539; // @[Mux.scala 31:69:@36574.4]
  assign _T_90541 = loadRequest_11 ? 16'h400 : _T_90540; // @[Mux.scala 31:69:@36575.4]
  assign _T_90542 = loadRequest_10 ? 16'h200 : _T_90541; // @[Mux.scala 31:69:@36576.4]
  assign _T_90543 = loadRequest_9 ? 16'h100 : _T_90542; // @[Mux.scala 31:69:@36577.4]
  assign _T_90544 = loadRequest_8 ? 16'h80 : _T_90543; // @[Mux.scala 31:69:@36578.4]
  assign _T_90545 = loadRequest_7 ? 16'h40 : _T_90544; // @[Mux.scala 31:69:@36579.4]
  assign _T_90546 = loadRequest_6 ? 16'h20 : _T_90545; // @[Mux.scala 31:69:@36580.4]
  assign _T_90547 = loadRequest_5 ? 16'h10 : _T_90546; // @[Mux.scala 31:69:@36581.4]
  assign _T_90548 = loadRequest_4 ? 16'h8 : _T_90547; // @[Mux.scala 31:69:@36582.4]
  assign _T_90549 = loadRequest_3 ? 16'h4 : _T_90548; // @[Mux.scala 31:69:@36583.4]
  assign _T_90550 = loadRequest_2 ? 16'h2 : _T_90549; // @[Mux.scala 31:69:@36584.4]
  assign _T_90551 = loadRequest_1 ? 16'h1 : _T_90550; // @[Mux.scala 31:69:@36585.4]
  assign _T_90552 = _T_90551[0]; // @[OneHot.scala 66:30:@36586.4]
  assign _T_90553 = _T_90551[1]; // @[OneHot.scala 66:30:@36587.4]
  assign _T_90554 = _T_90551[2]; // @[OneHot.scala 66:30:@36588.4]
  assign _T_90555 = _T_90551[3]; // @[OneHot.scala 66:30:@36589.4]
  assign _T_90556 = _T_90551[4]; // @[OneHot.scala 66:30:@36590.4]
  assign _T_90557 = _T_90551[5]; // @[OneHot.scala 66:30:@36591.4]
  assign _T_90558 = _T_90551[6]; // @[OneHot.scala 66:30:@36592.4]
  assign _T_90559 = _T_90551[7]; // @[OneHot.scala 66:30:@36593.4]
  assign _T_90560 = _T_90551[8]; // @[OneHot.scala 66:30:@36594.4]
  assign _T_90561 = _T_90551[9]; // @[OneHot.scala 66:30:@36595.4]
  assign _T_90562 = _T_90551[10]; // @[OneHot.scala 66:30:@36596.4]
  assign _T_90563 = _T_90551[11]; // @[OneHot.scala 66:30:@36597.4]
  assign _T_90564 = _T_90551[12]; // @[OneHot.scala 66:30:@36598.4]
  assign _T_90565 = _T_90551[13]; // @[OneHot.scala 66:30:@36599.4]
  assign _T_90566 = _T_90551[14]; // @[OneHot.scala 66:30:@36600.4]
  assign _T_90567 = _T_90551[15]; // @[OneHot.scala 66:30:@36601.4]
  assign _T_90608 = loadRequest_1 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36619.4]
  assign _T_90609 = loadRequest_0 ? 16'h4000 : _T_90608; // @[Mux.scala 31:69:@36620.4]
  assign _T_90610 = loadRequest_15 ? 16'h2000 : _T_90609; // @[Mux.scala 31:69:@36621.4]
  assign _T_90611 = loadRequest_14 ? 16'h1000 : _T_90610; // @[Mux.scala 31:69:@36622.4]
  assign _T_90612 = loadRequest_13 ? 16'h800 : _T_90611; // @[Mux.scala 31:69:@36623.4]
  assign _T_90613 = loadRequest_12 ? 16'h400 : _T_90612; // @[Mux.scala 31:69:@36624.4]
  assign _T_90614 = loadRequest_11 ? 16'h200 : _T_90613; // @[Mux.scala 31:69:@36625.4]
  assign _T_90615 = loadRequest_10 ? 16'h100 : _T_90614; // @[Mux.scala 31:69:@36626.4]
  assign _T_90616 = loadRequest_9 ? 16'h80 : _T_90615; // @[Mux.scala 31:69:@36627.4]
  assign _T_90617 = loadRequest_8 ? 16'h40 : _T_90616; // @[Mux.scala 31:69:@36628.4]
  assign _T_90618 = loadRequest_7 ? 16'h20 : _T_90617; // @[Mux.scala 31:69:@36629.4]
  assign _T_90619 = loadRequest_6 ? 16'h10 : _T_90618; // @[Mux.scala 31:69:@36630.4]
  assign _T_90620 = loadRequest_5 ? 16'h8 : _T_90619; // @[Mux.scala 31:69:@36631.4]
  assign _T_90621 = loadRequest_4 ? 16'h4 : _T_90620; // @[Mux.scala 31:69:@36632.4]
  assign _T_90622 = loadRequest_3 ? 16'h2 : _T_90621; // @[Mux.scala 31:69:@36633.4]
  assign _T_90623 = loadRequest_2 ? 16'h1 : _T_90622; // @[Mux.scala 31:69:@36634.4]
  assign _T_90624 = _T_90623[0]; // @[OneHot.scala 66:30:@36635.4]
  assign _T_90625 = _T_90623[1]; // @[OneHot.scala 66:30:@36636.4]
  assign _T_90626 = _T_90623[2]; // @[OneHot.scala 66:30:@36637.4]
  assign _T_90627 = _T_90623[3]; // @[OneHot.scala 66:30:@36638.4]
  assign _T_90628 = _T_90623[4]; // @[OneHot.scala 66:30:@36639.4]
  assign _T_90629 = _T_90623[5]; // @[OneHot.scala 66:30:@36640.4]
  assign _T_90630 = _T_90623[6]; // @[OneHot.scala 66:30:@36641.4]
  assign _T_90631 = _T_90623[7]; // @[OneHot.scala 66:30:@36642.4]
  assign _T_90632 = _T_90623[8]; // @[OneHot.scala 66:30:@36643.4]
  assign _T_90633 = _T_90623[9]; // @[OneHot.scala 66:30:@36644.4]
  assign _T_90634 = _T_90623[10]; // @[OneHot.scala 66:30:@36645.4]
  assign _T_90635 = _T_90623[11]; // @[OneHot.scala 66:30:@36646.4]
  assign _T_90636 = _T_90623[12]; // @[OneHot.scala 66:30:@36647.4]
  assign _T_90637 = _T_90623[13]; // @[OneHot.scala 66:30:@36648.4]
  assign _T_90638 = _T_90623[14]; // @[OneHot.scala 66:30:@36649.4]
  assign _T_90639 = _T_90623[15]; // @[OneHot.scala 66:30:@36650.4]
  assign _T_90680 = loadRequest_2 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36668.4]
  assign _T_90681 = loadRequest_1 ? 16'h4000 : _T_90680; // @[Mux.scala 31:69:@36669.4]
  assign _T_90682 = loadRequest_0 ? 16'h2000 : _T_90681; // @[Mux.scala 31:69:@36670.4]
  assign _T_90683 = loadRequest_15 ? 16'h1000 : _T_90682; // @[Mux.scala 31:69:@36671.4]
  assign _T_90684 = loadRequest_14 ? 16'h800 : _T_90683; // @[Mux.scala 31:69:@36672.4]
  assign _T_90685 = loadRequest_13 ? 16'h400 : _T_90684; // @[Mux.scala 31:69:@36673.4]
  assign _T_90686 = loadRequest_12 ? 16'h200 : _T_90685; // @[Mux.scala 31:69:@36674.4]
  assign _T_90687 = loadRequest_11 ? 16'h100 : _T_90686; // @[Mux.scala 31:69:@36675.4]
  assign _T_90688 = loadRequest_10 ? 16'h80 : _T_90687; // @[Mux.scala 31:69:@36676.4]
  assign _T_90689 = loadRequest_9 ? 16'h40 : _T_90688; // @[Mux.scala 31:69:@36677.4]
  assign _T_90690 = loadRequest_8 ? 16'h20 : _T_90689; // @[Mux.scala 31:69:@36678.4]
  assign _T_90691 = loadRequest_7 ? 16'h10 : _T_90690; // @[Mux.scala 31:69:@36679.4]
  assign _T_90692 = loadRequest_6 ? 16'h8 : _T_90691; // @[Mux.scala 31:69:@36680.4]
  assign _T_90693 = loadRequest_5 ? 16'h4 : _T_90692; // @[Mux.scala 31:69:@36681.4]
  assign _T_90694 = loadRequest_4 ? 16'h2 : _T_90693; // @[Mux.scala 31:69:@36682.4]
  assign _T_90695 = loadRequest_3 ? 16'h1 : _T_90694; // @[Mux.scala 31:69:@36683.4]
  assign _T_90696 = _T_90695[0]; // @[OneHot.scala 66:30:@36684.4]
  assign _T_90697 = _T_90695[1]; // @[OneHot.scala 66:30:@36685.4]
  assign _T_90698 = _T_90695[2]; // @[OneHot.scala 66:30:@36686.4]
  assign _T_90699 = _T_90695[3]; // @[OneHot.scala 66:30:@36687.4]
  assign _T_90700 = _T_90695[4]; // @[OneHot.scala 66:30:@36688.4]
  assign _T_90701 = _T_90695[5]; // @[OneHot.scala 66:30:@36689.4]
  assign _T_90702 = _T_90695[6]; // @[OneHot.scala 66:30:@36690.4]
  assign _T_90703 = _T_90695[7]; // @[OneHot.scala 66:30:@36691.4]
  assign _T_90704 = _T_90695[8]; // @[OneHot.scala 66:30:@36692.4]
  assign _T_90705 = _T_90695[9]; // @[OneHot.scala 66:30:@36693.4]
  assign _T_90706 = _T_90695[10]; // @[OneHot.scala 66:30:@36694.4]
  assign _T_90707 = _T_90695[11]; // @[OneHot.scala 66:30:@36695.4]
  assign _T_90708 = _T_90695[12]; // @[OneHot.scala 66:30:@36696.4]
  assign _T_90709 = _T_90695[13]; // @[OneHot.scala 66:30:@36697.4]
  assign _T_90710 = _T_90695[14]; // @[OneHot.scala 66:30:@36698.4]
  assign _T_90711 = _T_90695[15]; // @[OneHot.scala 66:30:@36699.4]
  assign _T_90752 = loadRequest_3 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36717.4]
  assign _T_90753 = loadRequest_2 ? 16'h4000 : _T_90752; // @[Mux.scala 31:69:@36718.4]
  assign _T_90754 = loadRequest_1 ? 16'h2000 : _T_90753; // @[Mux.scala 31:69:@36719.4]
  assign _T_90755 = loadRequest_0 ? 16'h1000 : _T_90754; // @[Mux.scala 31:69:@36720.4]
  assign _T_90756 = loadRequest_15 ? 16'h800 : _T_90755; // @[Mux.scala 31:69:@36721.4]
  assign _T_90757 = loadRequest_14 ? 16'h400 : _T_90756; // @[Mux.scala 31:69:@36722.4]
  assign _T_90758 = loadRequest_13 ? 16'h200 : _T_90757; // @[Mux.scala 31:69:@36723.4]
  assign _T_90759 = loadRequest_12 ? 16'h100 : _T_90758; // @[Mux.scala 31:69:@36724.4]
  assign _T_90760 = loadRequest_11 ? 16'h80 : _T_90759; // @[Mux.scala 31:69:@36725.4]
  assign _T_90761 = loadRequest_10 ? 16'h40 : _T_90760; // @[Mux.scala 31:69:@36726.4]
  assign _T_90762 = loadRequest_9 ? 16'h20 : _T_90761; // @[Mux.scala 31:69:@36727.4]
  assign _T_90763 = loadRequest_8 ? 16'h10 : _T_90762; // @[Mux.scala 31:69:@36728.4]
  assign _T_90764 = loadRequest_7 ? 16'h8 : _T_90763; // @[Mux.scala 31:69:@36729.4]
  assign _T_90765 = loadRequest_6 ? 16'h4 : _T_90764; // @[Mux.scala 31:69:@36730.4]
  assign _T_90766 = loadRequest_5 ? 16'h2 : _T_90765; // @[Mux.scala 31:69:@36731.4]
  assign _T_90767 = loadRequest_4 ? 16'h1 : _T_90766; // @[Mux.scala 31:69:@36732.4]
  assign _T_90768 = _T_90767[0]; // @[OneHot.scala 66:30:@36733.4]
  assign _T_90769 = _T_90767[1]; // @[OneHot.scala 66:30:@36734.4]
  assign _T_90770 = _T_90767[2]; // @[OneHot.scala 66:30:@36735.4]
  assign _T_90771 = _T_90767[3]; // @[OneHot.scala 66:30:@36736.4]
  assign _T_90772 = _T_90767[4]; // @[OneHot.scala 66:30:@36737.4]
  assign _T_90773 = _T_90767[5]; // @[OneHot.scala 66:30:@36738.4]
  assign _T_90774 = _T_90767[6]; // @[OneHot.scala 66:30:@36739.4]
  assign _T_90775 = _T_90767[7]; // @[OneHot.scala 66:30:@36740.4]
  assign _T_90776 = _T_90767[8]; // @[OneHot.scala 66:30:@36741.4]
  assign _T_90777 = _T_90767[9]; // @[OneHot.scala 66:30:@36742.4]
  assign _T_90778 = _T_90767[10]; // @[OneHot.scala 66:30:@36743.4]
  assign _T_90779 = _T_90767[11]; // @[OneHot.scala 66:30:@36744.4]
  assign _T_90780 = _T_90767[12]; // @[OneHot.scala 66:30:@36745.4]
  assign _T_90781 = _T_90767[13]; // @[OneHot.scala 66:30:@36746.4]
  assign _T_90782 = _T_90767[14]; // @[OneHot.scala 66:30:@36747.4]
  assign _T_90783 = _T_90767[15]; // @[OneHot.scala 66:30:@36748.4]
  assign _T_90824 = loadRequest_4 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36766.4]
  assign _T_90825 = loadRequest_3 ? 16'h4000 : _T_90824; // @[Mux.scala 31:69:@36767.4]
  assign _T_90826 = loadRequest_2 ? 16'h2000 : _T_90825; // @[Mux.scala 31:69:@36768.4]
  assign _T_90827 = loadRequest_1 ? 16'h1000 : _T_90826; // @[Mux.scala 31:69:@36769.4]
  assign _T_90828 = loadRequest_0 ? 16'h800 : _T_90827; // @[Mux.scala 31:69:@36770.4]
  assign _T_90829 = loadRequest_15 ? 16'h400 : _T_90828; // @[Mux.scala 31:69:@36771.4]
  assign _T_90830 = loadRequest_14 ? 16'h200 : _T_90829; // @[Mux.scala 31:69:@36772.4]
  assign _T_90831 = loadRequest_13 ? 16'h100 : _T_90830; // @[Mux.scala 31:69:@36773.4]
  assign _T_90832 = loadRequest_12 ? 16'h80 : _T_90831; // @[Mux.scala 31:69:@36774.4]
  assign _T_90833 = loadRequest_11 ? 16'h40 : _T_90832; // @[Mux.scala 31:69:@36775.4]
  assign _T_90834 = loadRequest_10 ? 16'h20 : _T_90833; // @[Mux.scala 31:69:@36776.4]
  assign _T_90835 = loadRequest_9 ? 16'h10 : _T_90834; // @[Mux.scala 31:69:@36777.4]
  assign _T_90836 = loadRequest_8 ? 16'h8 : _T_90835; // @[Mux.scala 31:69:@36778.4]
  assign _T_90837 = loadRequest_7 ? 16'h4 : _T_90836; // @[Mux.scala 31:69:@36779.4]
  assign _T_90838 = loadRequest_6 ? 16'h2 : _T_90837; // @[Mux.scala 31:69:@36780.4]
  assign _T_90839 = loadRequest_5 ? 16'h1 : _T_90838; // @[Mux.scala 31:69:@36781.4]
  assign _T_90840 = _T_90839[0]; // @[OneHot.scala 66:30:@36782.4]
  assign _T_90841 = _T_90839[1]; // @[OneHot.scala 66:30:@36783.4]
  assign _T_90842 = _T_90839[2]; // @[OneHot.scala 66:30:@36784.4]
  assign _T_90843 = _T_90839[3]; // @[OneHot.scala 66:30:@36785.4]
  assign _T_90844 = _T_90839[4]; // @[OneHot.scala 66:30:@36786.4]
  assign _T_90845 = _T_90839[5]; // @[OneHot.scala 66:30:@36787.4]
  assign _T_90846 = _T_90839[6]; // @[OneHot.scala 66:30:@36788.4]
  assign _T_90847 = _T_90839[7]; // @[OneHot.scala 66:30:@36789.4]
  assign _T_90848 = _T_90839[8]; // @[OneHot.scala 66:30:@36790.4]
  assign _T_90849 = _T_90839[9]; // @[OneHot.scala 66:30:@36791.4]
  assign _T_90850 = _T_90839[10]; // @[OneHot.scala 66:30:@36792.4]
  assign _T_90851 = _T_90839[11]; // @[OneHot.scala 66:30:@36793.4]
  assign _T_90852 = _T_90839[12]; // @[OneHot.scala 66:30:@36794.4]
  assign _T_90853 = _T_90839[13]; // @[OneHot.scala 66:30:@36795.4]
  assign _T_90854 = _T_90839[14]; // @[OneHot.scala 66:30:@36796.4]
  assign _T_90855 = _T_90839[15]; // @[OneHot.scala 66:30:@36797.4]
  assign _T_90896 = loadRequest_5 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36815.4]
  assign _T_90897 = loadRequest_4 ? 16'h4000 : _T_90896; // @[Mux.scala 31:69:@36816.4]
  assign _T_90898 = loadRequest_3 ? 16'h2000 : _T_90897; // @[Mux.scala 31:69:@36817.4]
  assign _T_90899 = loadRequest_2 ? 16'h1000 : _T_90898; // @[Mux.scala 31:69:@36818.4]
  assign _T_90900 = loadRequest_1 ? 16'h800 : _T_90899; // @[Mux.scala 31:69:@36819.4]
  assign _T_90901 = loadRequest_0 ? 16'h400 : _T_90900; // @[Mux.scala 31:69:@36820.4]
  assign _T_90902 = loadRequest_15 ? 16'h200 : _T_90901; // @[Mux.scala 31:69:@36821.4]
  assign _T_90903 = loadRequest_14 ? 16'h100 : _T_90902; // @[Mux.scala 31:69:@36822.4]
  assign _T_90904 = loadRequest_13 ? 16'h80 : _T_90903; // @[Mux.scala 31:69:@36823.4]
  assign _T_90905 = loadRequest_12 ? 16'h40 : _T_90904; // @[Mux.scala 31:69:@36824.4]
  assign _T_90906 = loadRequest_11 ? 16'h20 : _T_90905; // @[Mux.scala 31:69:@36825.4]
  assign _T_90907 = loadRequest_10 ? 16'h10 : _T_90906; // @[Mux.scala 31:69:@36826.4]
  assign _T_90908 = loadRequest_9 ? 16'h8 : _T_90907; // @[Mux.scala 31:69:@36827.4]
  assign _T_90909 = loadRequest_8 ? 16'h4 : _T_90908; // @[Mux.scala 31:69:@36828.4]
  assign _T_90910 = loadRequest_7 ? 16'h2 : _T_90909; // @[Mux.scala 31:69:@36829.4]
  assign _T_90911 = loadRequest_6 ? 16'h1 : _T_90910; // @[Mux.scala 31:69:@36830.4]
  assign _T_90912 = _T_90911[0]; // @[OneHot.scala 66:30:@36831.4]
  assign _T_90913 = _T_90911[1]; // @[OneHot.scala 66:30:@36832.4]
  assign _T_90914 = _T_90911[2]; // @[OneHot.scala 66:30:@36833.4]
  assign _T_90915 = _T_90911[3]; // @[OneHot.scala 66:30:@36834.4]
  assign _T_90916 = _T_90911[4]; // @[OneHot.scala 66:30:@36835.4]
  assign _T_90917 = _T_90911[5]; // @[OneHot.scala 66:30:@36836.4]
  assign _T_90918 = _T_90911[6]; // @[OneHot.scala 66:30:@36837.4]
  assign _T_90919 = _T_90911[7]; // @[OneHot.scala 66:30:@36838.4]
  assign _T_90920 = _T_90911[8]; // @[OneHot.scala 66:30:@36839.4]
  assign _T_90921 = _T_90911[9]; // @[OneHot.scala 66:30:@36840.4]
  assign _T_90922 = _T_90911[10]; // @[OneHot.scala 66:30:@36841.4]
  assign _T_90923 = _T_90911[11]; // @[OneHot.scala 66:30:@36842.4]
  assign _T_90924 = _T_90911[12]; // @[OneHot.scala 66:30:@36843.4]
  assign _T_90925 = _T_90911[13]; // @[OneHot.scala 66:30:@36844.4]
  assign _T_90926 = _T_90911[14]; // @[OneHot.scala 66:30:@36845.4]
  assign _T_90927 = _T_90911[15]; // @[OneHot.scala 66:30:@36846.4]
  assign _T_90968 = loadRequest_6 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36864.4]
  assign _T_90969 = loadRequest_5 ? 16'h4000 : _T_90968; // @[Mux.scala 31:69:@36865.4]
  assign _T_90970 = loadRequest_4 ? 16'h2000 : _T_90969; // @[Mux.scala 31:69:@36866.4]
  assign _T_90971 = loadRequest_3 ? 16'h1000 : _T_90970; // @[Mux.scala 31:69:@36867.4]
  assign _T_90972 = loadRequest_2 ? 16'h800 : _T_90971; // @[Mux.scala 31:69:@36868.4]
  assign _T_90973 = loadRequest_1 ? 16'h400 : _T_90972; // @[Mux.scala 31:69:@36869.4]
  assign _T_90974 = loadRequest_0 ? 16'h200 : _T_90973; // @[Mux.scala 31:69:@36870.4]
  assign _T_90975 = loadRequest_15 ? 16'h100 : _T_90974; // @[Mux.scala 31:69:@36871.4]
  assign _T_90976 = loadRequest_14 ? 16'h80 : _T_90975; // @[Mux.scala 31:69:@36872.4]
  assign _T_90977 = loadRequest_13 ? 16'h40 : _T_90976; // @[Mux.scala 31:69:@36873.4]
  assign _T_90978 = loadRequest_12 ? 16'h20 : _T_90977; // @[Mux.scala 31:69:@36874.4]
  assign _T_90979 = loadRequest_11 ? 16'h10 : _T_90978; // @[Mux.scala 31:69:@36875.4]
  assign _T_90980 = loadRequest_10 ? 16'h8 : _T_90979; // @[Mux.scala 31:69:@36876.4]
  assign _T_90981 = loadRequest_9 ? 16'h4 : _T_90980; // @[Mux.scala 31:69:@36877.4]
  assign _T_90982 = loadRequest_8 ? 16'h2 : _T_90981; // @[Mux.scala 31:69:@36878.4]
  assign _T_90983 = loadRequest_7 ? 16'h1 : _T_90982; // @[Mux.scala 31:69:@36879.4]
  assign _T_90984 = _T_90983[0]; // @[OneHot.scala 66:30:@36880.4]
  assign _T_90985 = _T_90983[1]; // @[OneHot.scala 66:30:@36881.4]
  assign _T_90986 = _T_90983[2]; // @[OneHot.scala 66:30:@36882.4]
  assign _T_90987 = _T_90983[3]; // @[OneHot.scala 66:30:@36883.4]
  assign _T_90988 = _T_90983[4]; // @[OneHot.scala 66:30:@36884.4]
  assign _T_90989 = _T_90983[5]; // @[OneHot.scala 66:30:@36885.4]
  assign _T_90990 = _T_90983[6]; // @[OneHot.scala 66:30:@36886.4]
  assign _T_90991 = _T_90983[7]; // @[OneHot.scala 66:30:@36887.4]
  assign _T_90992 = _T_90983[8]; // @[OneHot.scala 66:30:@36888.4]
  assign _T_90993 = _T_90983[9]; // @[OneHot.scala 66:30:@36889.4]
  assign _T_90994 = _T_90983[10]; // @[OneHot.scala 66:30:@36890.4]
  assign _T_90995 = _T_90983[11]; // @[OneHot.scala 66:30:@36891.4]
  assign _T_90996 = _T_90983[12]; // @[OneHot.scala 66:30:@36892.4]
  assign _T_90997 = _T_90983[13]; // @[OneHot.scala 66:30:@36893.4]
  assign _T_90998 = _T_90983[14]; // @[OneHot.scala 66:30:@36894.4]
  assign _T_90999 = _T_90983[15]; // @[OneHot.scala 66:30:@36895.4]
  assign _T_91040 = loadRequest_7 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36913.4]
  assign _T_91041 = loadRequest_6 ? 16'h4000 : _T_91040; // @[Mux.scala 31:69:@36914.4]
  assign _T_91042 = loadRequest_5 ? 16'h2000 : _T_91041; // @[Mux.scala 31:69:@36915.4]
  assign _T_91043 = loadRequest_4 ? 16'h1000 : _T_91042; // @[Mux.scala 31:69:@36916.4]
  assign _T_91044 = loadRequest_3 ? 16'h800 : _T_91043; // @[Mux.scala 31:69:@36917.4]
  assign _T_91045 = loadRequest_2 ? 16'h400 : _T_91044; // @[Mux.scala 31:69:@36918.4]
  assign _T_91046 = loadRequest_1 ? 16'h200 : _T_91045; // @[Mux.scala 31:69:@36919.4]
  assign _T_91047 = loadRequest_0 ? 16'h100 : _T_91046; // @[Mux.scala 31:69:@36920.4]
  assign _T_91048 = loadRequest_15 ? 16'h80 : _T_91047; // @[Mux.scala 31:69:@36921.4]
  assign _T_91049 = loadRequest_14 ? 16'h40 : _T_91048; // @[Mux.scala 31:69:@36922.4]
  assign _T_91050 = loadRequest_13 ? 16'h20 : _T_91049; // @[Mux.scala 31:69:@36923.4]
  assign _T_91051 = loadRequest_12 ? 16'h10 : _T_91050; // @[Mux.scala 31:69:@36924.4]
  assign _T_91052 = loadRequest_11 ? 16'h8 : _T_91051; // @[Mux.scala 31:69:@36925.4]
  assign _T_91053 = loadRequest_10 ? 16'h4 : _T_91052; // @[Mux.scala 31:69:@36926.4]
  assign _T_91054 = loadRequest_9 ? 16'h2 : _T_91053; // @[Mux.scala 31:69:@36927.4]
  assign _T_91055 = loadRequest_8 ? 16'h1 : _T_91054; // @[Mux.scala 31:69:@36928.4]
  assign _T_91056 = _T_91055[0]; // @[OneHot.scala 66:30:@36929.4]
  assign _T_91057 = _T_91055[1]; // @[OneHot.scala 66:30:@36930.4]
  assign _T_91058 = _T_91055[2]; // @[OneHot.scala 66:30:@36931.4]
  assign _T_91059 = _T_91055[3]; // @[OneHot.scala 66:30:@36932.4]
  assign _T_91060 = _T_91055[4]; // @[OneHot.scala 66:30:@36933.4]
  assign _T_91061 = _T_91055[5]; // @[OneHot.scala 66:30:@36934.4]
  assign _T_91062 = _T_91055[6]; // @[OneHot.scala 66:30:@36935.4]
  assign _T_91063 = _T_91055[7]; // @[OneHot.scala 66:30:@36936.4]
  assign _T_91064 = _T_91055[8]; // @[OneHot.scala 66:30:@36937.4]
  assign _T_91065 = _T_91055[9]; // @[OneHot.scala 66:30:@36938.4]
  assign _T_91066 = _T_91055[10]; // @[OneHot.scala 66:30:@36939.4]
  assign _T_91067 = _T_91055[11]; // @[OneHot.scala 66:30:@36940.4]
  assign _T_91068 = _T_91055[12]; // @[OneHot.scala 66:30:@36941.4]
  assign _T_91069 = _T_91055[13]; // @[OneHot.scala 66:30:@36942.4]
  assign _T_91070 = _T_91055[14]; // @[OneHot.scala 66:30:@36943.4]
  assign _T_91071 = _T_91055[15]; // @[OneHot.scala 66:30:@36944.4]
  assign _T_91112 = loadRequest_8 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36962.4]
  assign _T_91113 = loadRequest_7 ? 16'h4000 : _T_91112; // @[Mux.scala 31:69:@36963.4]
  assign _T_91114 = loadRequest_6 ? 16'h2000 : _T_91113; // @[Mux.scala 31:69:@36964.4]
  assign _T_91115 = loadRequest_5 ? 16'h1000 : _T_91114; // @[Mux.scala 31:69:@36965.4]
  assign _T_91116 = loadRequest_4 ? 16'h800 : _T_91115; // @[Mux.scala 31:69:@36966.4]
  assign _T_91117 = loadRequest_3 ? 16'h400 : _T_91116; // @[Mux.scala 31:69:@36967.4]
  assign _T_91118 = loadRequest_2 ? 16'h200 : _T_91117; // @[Mux.scala 31:69:@36968.4]
  assign _T_91119 = loadRequest_1 ? 16'h100 : _T_91118; // @[Mux.scala 31:69:@36969.4]
  assign _T_91120 = loadRequest_0 ? 16'h80 : _T_91119; // @[Mux.scala 31:69:@36970.4]
  assign _T_91121 = loadRequest_15 ? 16'h40 : _T_91120; // @[Mux.scala 31:69:@36971.4]
  assign _T_91122 = loadRequest_14 ? 16'h20 : _T_91121; // @[Mux.scala 31:69:@36972.4]
  assign _T_91123 = loadRequest_13 ? 16'h10 : _T_91122; // @[Mux.scala 31:69:@36973.4]
  assign _T_91124 = loadRequest_12 ? 16'h8 : _T_91123; // @[Mux.scala 31:69:@36974.4]
  assign _T_91125 = loadRequest_11 ? 16'h4 : _T_91124; // @[Mux.scala 31:69:@36975.4]
  assign _T_91126 = loadRequest_10 ? 16'h2 : _T_91125; // @[Mux.scala 31:69:@36976.4]
  assign _T_91127 = loadRequest_9 ? 16'h1 : _T_91126; // @[Mux.scala 31:69:@36977.4]
  assign _T_91128 = _T_91127[0]; // @[OneHot.scala 66:30:@36978.4]
  assign _T_91129 = _T_91127[1]; // @[OneHot.scala 66:30:@36979.4]
  assign _T_91130 = _T_91127[2]; // @[OneHot.scala 66:30:@36980.4]
  assign _T_91131 = _T_91127[3]; // @[OneHot.scala 66:30:@36981.4]
  assign _T_91132 = _T_91127[4]; // @[OneHot.scala 66:30:@36982.4]
  assign _T_91133 = _T_91127[5]; // @[OneHot.scala 66:30:@36983.4]
  assign _T_91134 = _T_91127[6]; // @[OneHot.scala 66:30:@36984.4]
  assign _T_91135 = _T_91127[7]; // @[OneHot.scala 66:30:@36985.4]
  assign _T_91136 = _T_91127[8]; // @[OneHot.scala 66:30:@36986.4]
  assign _T_91137 = _T_91127[9]; // @[OneHot.scala 66:30:@36987.4]
  assign _T_91138 = _T_91127[10]; // @[OneHot.scala 66:30:@36988.4]
  assign _T_91139 = _T_91127[11]; // @[OneHot.scala 66:30:@36989.4]
  assign _T_91140 = _T_91127[12]; // @[OneHot.scala 66:30:@36990.4]
  assign _T_91141 = _T_91127[13]; // @[OneHot.scala 66:30:@36991.4]
  assign _T_91142 = _T_91127[14]; // @[OneHot.scala 66:30:@36992.4]
  assign _T_91143 = _T_91127[15]; // @[OneHot.scala 66:30:@36993.4]
  assign _T_91184 = loadRequest_9 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37011.4]
  assign _T_91185 = loadRequest_8 ? 16'h4000 : _T_91184; // @[Mux.scala 31:69:@37012.4]
  assign _T_91186 = loadRequest_7 ? 16'h2000 : _T_91185; // @[Mux.scala 31:69:@37013.4]
  assign _T_91187 = loadRequest_6 ? 16'h1000 : _T_91186; // @[Mux.scala 31:69:@37014.4]
  assign _T_91188 = loadRequest_5 ? 16'h800 : _T_91187; // @[Mux.scala 31:69:@37015.4]
  assign _T_91189 = loadRequest_4 ? 16'h400 : _T_91188; // @[Mux.scala 31:69:@37016.4]
  assign _T_91190 = loadRequest_3 ? 16'h200 : _T_91189; // @[Mux.scala 31:69:@37017.4]
  assign _T_91191 = loadRequest_2 ? 16'h100 : _T_91190; // @[Mux.scala 31:69:@37018.4]
  assign _T_91192 = loadRequest_1 ? 16'h80 : _T_91191; // @[Mux.scala 31:69:@37019.4]
  assign _T_91193 = loadRequest_0 ? 16'h40 : _T_91192; // @[Mux.scala 31:69:@37020.4]
  assign _T_91194 = loadRequest_15 ? 16'h20 : _T_91193; // @[Mux.scala 31:69:@37021.4]
  assign _T_91195 = loadRequest_14 ? 16'h10 : _T_91194; // @[Mux.scala 31:69:@37022.4]
  assign _T_91196 = loadRequest_13 ? 16'h8 : _T_91195; // @[Mux.scala 31:69:@37023.4]
  assign _T_91197 = loadRequest_12 ? 16'h4 : _T_91196; // @[Mux.scala 31:69:@37024.4]
  assign _T_91198 = loadRequest_11 ? 16'h2 : _T_91197; // @[Mux.scala 31:69:@37025.4]
  assign _T_91199 = loadRequest_10 ? 16'h1 : _T_91198; // @[Mux.scala 31:69:@37026.4]
  assign _T_91200 = _T_91199[0]; // @[OneHot.scala 66:30:@37027.4]
  assign _T_91201 = _T_91199[1]; // @[OneHot.scala 66:30:@37028.4]
  assign _T_91202 = _T_91199[2]; // @[OneHot.scala 66:30:@37029.4]
  assign _T_91203 = _T_91199[3]; // @[OneHot.scala 66:30:@37030.4]
  assign _T_91204 = _T_91199[4]; // @[OneHot.scala 66:30:@37031.4]
  assign _T_91205 = _T_91199[5]; // @[OneHot.scala 66:30:@37032.4]
  assign _T_91206 = _T_91199[6]; // @[OneHot.scala 66:30:@37033.4]
  assign _T_91207 = _T_91199[7]; // @[OneHot.scala 66:30:@37034.4]
  assign _T_91208 = _T_91199[8]; // @[OneHot.scala 66:30:@37035.4]
  assign _T_91209 = _T_91199[9]; // @[OneHot.scala 66:30:@37036.4]
  assign _T_91210 = _T_91199[10]; // @[OneHot.scala 66:30:@37037.4]
  assign _T_91211 = _T_91199[11]; // @[OneHot.scala 66:30:@37038.4]
  assign _T_91212 = _T_91199[12]; // @[OneHot.scala 66:30:@37039.4]
  assign _T_91213 = _T_91199[13]; // @[OneHot.scala 66:30:@37040.4]
  assign _T_91214 = _T_91199[14]; // @[OneHot.scala 66:30:@37041.4]
  assign _T_91215 = _T_91199[15]; // @[OneHot.scala 66:30:@37042.4]
  assign _T_91256 = loadRequest_10 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37060.4]
  assign _T_91257 = loadRequest_9 ? 16'h4000 : _T_91256; // @[Mux.scala 31:69:@37061.4]
  assign _T_91258 = loadRequest_8 ? 16'h2000 : _T_91257; // @[Mux.scala 31:69:@37062.4]
  assign _T_91259 = loadRequest_7 ? 16'h1000 : _T_91258; // @[Mux.scala 31:69:@37063.4]
  assign _T_91260 = loadRequest_6 ? 16'h800 : _T_91259; // @[Mux.scala 31:69:@37064.4]
  assign _T_91261 = loadRequest_5 ? 16'h400 : _T_91260; // @[Mux.scala 31:69:@37065.4]
  assign _T_91262 = loadRequest_4 ? 16'h200 : _T_91261; // @[Mux.scala 31:69:@37066.4]
  assign _T_91263 = loadRequest_3 ? 16'h100 : _T_91262; // @[Mux.scala 31:69:@37067.4]
  assign _T_91264 = loadRequest_2 ? 16'h80 : _T_91263; // @[Mux.scala 31:69:@37068.4]
  assign _T_91265 = loadRequest_1 ? 16'h40 : _T_91264; // @[Mux.scala 31:69:@37069.4]
  assign _T_91266 = loadRequest_0 ? 16'h20 : _T_91265; // @[Mux.scala 31:69:@37070.4]
  assign _T_91267 = loadRequest_15 ? 16'h10 : _T_91266; // @[Mux.scala 31:69:@37071.4]
  assign _T_91268 = loadRequest_14 ? 16'h8 : _T_91267; // @[Mux.scala 31:69:@37072.4]
  assign _T_91269 = loadRequest_13 ? 16'h4 : _T_91268; // @[Mux.scala 31:69:@37073.4]
  assign _T_91270 = loadRequest_12 ? 16'h2 : _T_91269; // @[Mux.scala 31:69:@37074.4]
  assign _T_91271 = loadRequest_11 ? 16'h1 : _T_91270; // @[Mux.scala 31:69:@37075.4]
  assign _T_91272 = _T_91271[0]; // @[OneHot.scala 66:30:@37076.4]
  assign _T_91273 = _T_91271[1]; // @[OneHot.scala 66:30:@37077.4]
  assign _T_91274 = _T_91271[2]; // @[OneHot.scala 66:30:@37078.4]
  assign _T_91275 = _T_91271[3]; // @[OneHot.scala 66:30:@37079.4]
  assign _T_91276 = _T_91271[4]; // @[OneHot.scala 66:30:@37080.4]
  assign _T_91277 = _T_91271[5]; // @[OneHot.scala 66:30:@37081.4]
  assign _T_91278 = _T_91271[6]; // @[OneHot.scala 66:30:@37082.4]
  assign _T_91279 = _T_91271[7]; // @[OneHot.scala 66:30:@37083.4]
  assign _T_91280 = _T_91271[8]; // @[OneHot.scala 66:30:@37084.4]
  assign _T_91281 = _T_91271[9]; // @[OneHot.scala 66:30:@37085.4]
  assign _T_91282 = _T_91271[10]; // @[OneHot.scala 66:30:@37086.4]
  assign _T_91283 = _T_91271[11]; // @[OneHot.scala 66:30:@37087.4]
  assign _T_91284 = _T_91271[12]; // @[OneHot.scala 66:30:@37088.4]
  assign _T_91285 = _T_91271[13]; // @[OneHot.scala 66:30:@37089.4]
  assign _T_91286 = _T_91271[14]; // @[OneHot.scala 66:30:@37090.4]
  assign _T_91287 = _T_91271[15]; // @[OneHot.scala 66:30:@37091.4]
  assign _T_91328 = loadRequest_11 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37109.4]
  assign _T_91329 = loadRequest_10 ? 16'h4000 : _T_91328; // @[Mux.scala 31:69:@37110.4]
  assign _T_91330 = loadRequest_9 ? 16'h2000 : _T_91329; // @[Mux.scala 31:69:@37111.4]
  assign _T_91331 = loadRequest_8 ? 16'h1000 : _T_91330; // @[Mux.scala 31:69:@37112.4]
  assign _T_91332 = loadRequest_7 ? 16'h800 : _T_91331; // @[Mux.scala 31:69:@37113.4]
  assign _T_91333 = loadRequest_6 ? 16'h400 : _T_91332; // @[Mux.scala 31:69:@37114.4]
  assign _T_91334 = loadRequest_5 ? 16'h200 : _T_91333; // @[Mux.scala 31:69:@37115.4]
  assign _T_91335 = loadRequest_4 ? 16'h100 : _T_91334; // @[Mux.scala 31:69:@37116.4]
  assign _T_91336 = loadRequest_3 ? 16'h80 : _T_91335; // @[Mux.scala 31:69:@37117.4]
  assign _T_91337 = loadRequest_2 ? 16'h40 : _T_91336; // @[Mux.scala 31:69:@37118.4]
  assign _T_91338 = loadRequest_1 ? 16'h20 : _T_91337; // @[Mux.scala 31:69:@37119.4]
  assign _T_91339 = loadRequest_0 ? 16'h10 : _T_91338; // @[Mux.scala 31:69:@37120.4]
  assign _T_91340 = loadRequest_15 ? 16'h8 : _T_91339; // @[Mux.scala 31:69:@37121.4]
  assign _T_91341 = loadRequest_14 ? 16'h4 : _T_91340; // @[Mux.scala 31:69:@37122.4]
  assign _T_91342 = loadRequest_13 ? 16'h2 : _T_91341; // @[Mux.scala 31:69:@37123.4]
  assign _T_91343 = loadRequest_12 ? 16'h1 : _T_91342; // @[Mux.scala 31:69:@37124.4]
  assign _T_91344 = _T_91343[0]; // @[OneHot.scala 66:30:@37125.4]
  assign _T_91345 = _T_91343[1]; // @[OneHot.scala 66:30:@37126.4]
  assign _T_91346 = _T_91343[2]; // @[OneHot.scala 66:30:@37127.4]
  assign _T_91347 = _T_91343[3]; // @[OneHot.scala 66:30:@37128.4]
  assign _T_91348 = _T_91343[4]; // @[OneHot.scala 66:30:@37129.4]
  assign _T_91349 = _T_91343[5]; // @[OneHot.scala 66:30:@37130.4]
  assign _T_91350 = _T_91343[6]; // @[OneHot.scala 66:30:@37131.4]
  assign _T_91351 = _T_91343[7]; // @[OneHot.scala 66:30:@37132.4]
  assign _T_91352 = _T_91343[8]; // @[OneHot.scala 66:30:@37133.4]
  assign _T_91353 = _T_91343[9]; // @[OneHot.scala 66:30:@37134.4]
  assign _T_91354 = _T_91343[10]; // @[OneHot.scala 66:30:@37135.4]
  assign _T_91355 = _T_91343[11]; // @[OneHot.scala 66:30:@37136.4]
  assign _T_91356 = _T_91343[12]; // @[OneHot.scala 66:30:@37137.4]
  assign _T_91357 = _T_91343[13]; // @[OneHot.scala 66:30:@37138.4]
  assign _T_91358 = _T_91343[14]; // @[OneHot.scala 66:30:@37139.4]
  assign _T_91359 = _T_91343[15]; // @[OneHot.scala 66:30:@37140.4]
  assign _T_91400 = loadRequest_12 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37158.4]
  assign _T_91401 = loadRequest_11 ? 16'h4000 : _T_91400; // @[Mux.scala 31:69:@37159.4]
  assign _T_91402 = loadRequest_10 ? 16'h2000 : _T_91401; // @[Mux.scala 31:69:@37160.4]
  assign _T_91403 = loadRequest_9 ? 16'h1000 : _T_91402; // @[Mux.scala 31:69:@37161.4]
  assign _T_91404 = loadRequest_8 ? 16'h800 : _T_91403; // @[Mux.scala 31:69:@37162.4]
  assign _T_91405 = loadRequest_7 ? 16'h400 : _T_91404; // @[Mux.scala 31:69:@37163.4]
  assign _T_91406 = loadRequest_6 ? 16'h200 : _T_91405; // @[Mux.scala 31:69:@37164.4]
  assign _T_91407 = loadRequest_5 ? 16'h100 : _T_91406; // @[Mux.scala 31:69:@37165.4]
  assign _T_91408 = loadRequest_4 ? 16'h80 : _T_91407; // @[Mux.scala 31:69:@37166.4]
  assign _T_91409 = loadRequest_3 ? 16'h40 : _T_91408; // @[Mux.scala 31:69:@37167.4]
  assign _T_91410 = loadRequest_2 ? 16'h20 : _T_91409; // @[Mux.scala 31:69:@37168.4]
  assign _T_91411 = loadRequest_1 ? 16'h10 : _T_91410; // @[Mux.scala 31:69:@37169.4]
  assign _T_91412 = loadRequest_0 ? 16'h8 : _T_91411; // @[Mux.scala 31:69:@37170.4]
  assign _T_91413 = loadRequest_15 ? 16'h4 : _T_91412; // @[Mux.scala 31:69:@37171.4]
  assign _T_91414 = loadRequest_14 ? 16'h2 : _T_91413; // @[Mux.scala 31:69:@37172.4]
  assign _T_91415 = loadRequest_13 ? 16'h1 : _T_91414; // @[Mux.scala 31:69:@37173.4]
  assign _T_91416 = _T_91415[0]; // @[OneHot.scala 66:30:@37174.4]
  assign _T_91417 = _T_91415[1]; // @[OneHot.scala 66:30:@37175.4]
  assign _T_91418 = _T_91415[2]; // @[OneHot.scala 66:30:@37176.4]
  assign _T_91419 = _T_91415[3]; // @[OneHot.scala 66:30:@37177.4]
  assign _T_91420 = _T_91415[4]; // @[OneHot.scala 66:30:@37178.4]
  assign _T_91421 = _T_91415[5]; // @[OneHot.scala 66:30:@37179.4]
  assign _T_91422 = _T_91415[6]; // @[OneHot.scala 66:30:@37180.4]
  assign _T_91423 = _T_91415[7]; // @[OneHot.scala 66:30:@37181.4]
  assign _T_91424 = _T_91415[8]; // @[OneHot.scala 66:30:@37182.4]
  assign _T_91425 = _T_91415[9]; // @[OneHot.scala 66:30:@37183.4]
  assign _T_91426 = _T_91415[10]; // @[OneHot.scala 66:30:@37184.4]
  assign _T_91427 = _T_91415[11]; // @[OneHot.scala 66:30:@37185.4]
  assign _T_91428 = _T_91415[12]; // @[OneHot.scala 66:30:@37186.4]
  assign _T_91429 = _T_91415[13]; // @[OneHot.scala 66:30:@37187.4]
  assign _T_91430 = _T_91415[14]; // @[OneHot.scala 66:30:@37188.4]
  assign _T_91431 = _T_91415[15]; // @[OneHot.scala 66:30:@37189.4]
  assign _T_91472 = loadRequest_13 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37207.4]
  assign _T_91473 = loadRequest_12 ? 16'h4000 : _T_91472; // @[Mux.scala 31:69:@37208.4]
  assign _T_91474 = loadRequest_11 ? 16'h2000 : _T_91473; // @[Mux.scala 31:69:@37209.4]
  assign _T_91475 = loadRequest_10 ? 16'h1000 : _T_91474; // @[Mux.scala 31:69:@37210.4]
  assign _T_91476 = loadRequest_9 ? 16'h800 : _T_91475; // @[Mux.scala 31:69:@37211.4]
  assign _T_91477 = loadRequest_8 ? 16'h400 : _T_91476; // @[Mux.scala 31:69:@37212.4]
  assign _T_91478 = loadRequest_7 ? 16'h200 : _T_91477; // @[Mux.scala 31:69:@37213.4]
  assign _T_91479 = loadRequest_6 ? 16'h100 : _T_91478; // @[Mux.scala 31:69:@37214.4]
  assign _T_91480 = loadRequest_5 ? 16'h80 : _T_91479; // @[Mux.scala 31:69:@37215.4]
  assign _T_91481 = loadRequest_4 ? 16'h40 : _T_91480; // @[Mux.scala 31:69:@37216.4]
  assign _T_91482 = loadRequest_3 ? 16'h20 : _T_91481; // @[Mux.scala 31:69:@37217.4]
  assign _T_91483 = loadRequest_2 ? 16'h10 : _T_91482; // @[Mux.scala 31:69:@37218.4]
  assign _T_91484 = loadRequest_1 ? 16'h8 : _T_91483; // @[Mux.scala 31:69:@37219.4]
  assign _T_91485 = loadRequest_0 ? 16'h4 : _T_91484; // @[Mux.scala 31:69:@37220.4]
  assign _T_91486 = loadRequest_15 ? 16'h2 : _T_91485; // @[Mux.scala 31:69:@37221.4]
  assign _T_91487 = loadRequest_14 ? 16'h1 : _T_91486; // @[Mux.scala 31:69:@37222.4]
  assign _T_91488 = _T_91487[0]; // @[OneHot.scala 66:30:@37223.4]
  assign _T_91489 = _T_91487[1]; // @[OneHot.scala 66:30:@37224.4]
  assign _T_91490 = _T_91487[2]; // @[OneHot.scala 66:30:@37225.4]
  assign _T_91491 = _T_91487[3]; // @[OneHot.scala 66:30:@37226.4]
  assign _T_91492 = _T_91487[4]; // @[OneHot.scala 66:30:@37227.4]
  assign _T_91493 = _T_91487[5]; // @[OneHot.scala 66:30:@37228.4]
  assign _T_91494 = _T_91487[6]; // @[OneHot.scala 66:30:@37229.4]
  assign _T_91495 = _T_91487[7]; // @[OneHot.scala 66:30:@37230.4]
  assign _T_91496 = _T_91487[8]; // @[OneHot.scala 66:30:@37231.4]
  assign _T_91497 = _T_91487[9]; // @[OneHot.scala 66:30:@37232.4]
  assign _T_91498 = _T_91487[10]; // @[OneHot.scala 66:30:@37233.4]
  assign _T_91499 = _T_91487[11]; // @[OneHot.scala 66:30:@37234.4]
  assign _T_91500 = _T_91487[12]; // @[OneHot.scala 66:30:@37235.4]
  assign _T_91501 = _T_91487[13]; // @[OneHot.scala 66:30:@37236.4]
  assign _T_91502 = _T_91487[14]; // @[OneHot.scala 66:30:@37237.4]
  assign _T_91503 = _T_91487[15]; // @[OneHot.scala 66:30:@37238.4]
  assign _T_91544 = loadRequest_14 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37256.4]
  assign _T_91545 = loadRequest_13 ? 16'h4000 : _T_91544; // @[Mux.scala 31:69:@37257.4]
  assign _T_91546 = loadRequest_12 ? 16'h2000 : _T_91545; // @[Mux.scala 31:69:@37258.4]
  assign _T_91547 = loadRequest_11 ? 16'h1000 : _T_91546; // @[Mux.scala 31:69:@37259.4]
  assign _T_91548 = loadRequest_10 ? 16'h800 : _T_91547; // @[Mux.scala 31:69:@37260.4]
  assign _T_91549 = loadRequest_9 ? 16'h400 : _T_91548; // @[Mux.scala 31:69:@37261.4]
  assign _T_91550 = loadRequest_8 ? 16'h200 : _T_91549; // @[Mux.scala 31:69:@37262.4]
  assign _T_91551 = loadRequest_7 ? 16'h100 : _T_91550; // @[Mux.scala 31:69:@37263.4]
  assign _T_91552 = loadRequest_6 ? 16'h80 : _T_91551; // @[Mux.scala 31:69:@37264.4]
  assign _T_91553 = loadRequest_5 ? 16'h40 : _T_91552; // @[Mux.scala 31:69:@37265.4]
  assign _T_91554 = loadRequest_4 ? 16'h20 : _T_91553; // @[Mux.scala 31:69:@37266.4]
  assign _T_91555 = loadRequest_3 ? 16'h10 : _T_91554; // @[Mux.scala 31:69:@37267.4]
  assign _T_91556 = loadRequest_2 ? 16'h8 : _T_91555; // @[Mux.scala 31:69:@37268.4]
  assign _T_91557 = loadRequest_1 ? 16'h4 : _T_91556; // @[Mux.scala 31:69:@37269.4]
  assign _T_91558 = loadRequest_0 ? 16'h2 : _T_91557; // @[Mux.scala 31:69:@37270.4]
  assign _T_91559 = loadRequest_15 ? 16'h1 : _T_91558; // @[Mux.scala 31:69:@37271.4]
  assign _T_91560 = _T_91559[0]; // @[OneHot.scala 66:30:@37272.4]
  assign _T_91561 = _T_91559[1]; // @[OneHot.scala 66:30:@37273.4]
  assign _T_91562 = _T_91559[2]; // @[OneHot.scala 66:30:@37274.4]
  assign _T_91563 = _T_91559[3]; // @[OneHot.scala 66:30:@37275.4]
  assign _T_91564 = _T_91559[4]; // @[OneHot.scala 66:30:@37276.4]
  assign _T_91565 = _T_91559[5]; // @[OneHot.scala 66:30:@37277.4]
  assign _T_91566 = _T_91559[6]; // @[OneHot.scala 66:30:@37278.4]
  assign _T_91567 = _T_91559[7]; // @[OneHot.scala 66:30:@37279.4]
  assign _T_91568 = _T_91559[8]; // @[OneHot.scala 66:30:@37280.4]
  assign _T_91569 = _T_91559[9]; // @[OneHot.scala 66:30:@37281.4]
  assign _T_91570 = _T_91559[10]; // @[OneHot.scala 66:30:@37282.4]
  assign _T_91571 = _T_91559[11]; // @[OneHot.scala 66:30:@37283.4]
  assign _T_91572 = _T_91559[12]; // @[OneHot.scala 66:30:@37284.4]
  assign _T_91573 = _T_91559[13]; // @[OneHot.scala 66:30:@37285.4]
  assign _T_91574 = _T_91559[14]; // @[OneHot.scala 66:30:@37286.4]
  assign _T_91575 = _T_91559[15]; // @[OneHot.scala 66:30:@37287.4]
  assign _T_91640 = {_T_90487,_T_90486,_T_90485,_T_90484,_T_90483,_T_90482,_T_90481,_T_90480}; // @[Mux.scala 19:72:@37311.4]
  assign _T_91648 = {_T_90495,_T_90494,_T_90493,_T_90492,_T_90491,_T_90490,_T_90489,_T_90488,_T_91640}; // @[Mux.scala 19:72:@37319.4]
  assign _T_91650 = _T_90408 ? _T_91648 : 16'h0; // @[Mux.scala 19:72:@37320.4]
  assign _T_91657 = {_T_90558,_T_90557,_T_90556,_T_90555,_T_90554,_T_90553,_T_90552,_T_90567}; // @[Mux.scala 19:72:@37327.4]
  assign _T_91665 = {_T_90566,_T_90565,_T_90564,_T_90563,_T_90562,_T_90561,_T_90560,_T_90559,_T_91657}; // @[Mux.scala 19:72:@37335.4]
  assign _T_91667 = _T_90409 ? _T_91665 : 16'h0; // @[Mux.scala 19:72:@37336.4]
  assign _T_91674 = {_T_90629,_T_90628,_T_90627,_T_90626,_T_90625,_T_90624,_T_90639,_T_90638}; // @[Mux.scala 19:72:@37343.4]
  assign _T_91682 = {_T_90637,_T_90636,_T_90635,_T_90634,_T_90633,_T_90632,_T_90631,_T_90630,_T_91674}; // @[Mux.scala 19:72:@37351.4]
  assign _T_91684 = _T_90410 ? _T_91682 : 16'h0; // @[Mux.scala 19:72:@37352.4]
  assign _T_91691 = {_T_90700,_T_90699,_T_90698,_T_90697,_T_90696,_T_90711,_T_90710,_T_90709}; // @[Mux.scala 19:72:@37359.4]
  assign _T_91699 = {_T_90708,_T_90707,_T_90706,_T_90705,_T_90704,_T_90703,_T_90702,_T_90701,_T_91691}; // @[Mux.scala 19:72:@37367.4]
  assign _T_91701 = _T_90411 ? _T_91699 : 16'h0; // @[Mux.scala 19:72:@37368.4]
  assign _T_91708 = {_T_90771,_T_90770,_T_90769,_T_90768,_T_90783,_T_90782,_T_90781,_T_90780}; // @[Mux.scala 19:72:@37375.4]
  assign _T_91716 = {_T_90779,_T_90778,_T_90777,_T_90776,_T_90775,_T_90774,_T_90773,_T_90772,_T_91708}; // @[Mux.scala 19:72:@37383.4]
  assign _T_91718 = _T_90412 ? _T_91716 : 16'h0; // @[Mux.scala 19:72:@37384.4]
  assign _T_91725 = {_T_90842,_T_90841,_T_90840,_T_90855,_T_90854,_T_90853,_T_90852,_T_90851}; // @[Mux.scala 19:72:@37391.4]
  assign _T_91733 = {_T_90850,_T_90849,_T_90848,_T_90847,_T_90846,_T_90845,_T_90844,_T_90843,_T_91725}; // @[Mux.scala 19:72:@37399.4]
  assign _T_91735 = _T_90413 ? _T_91733 : 16'h0; // @[Mux.scala 19:72:@37400.4]
  assign _T_91742 = {_T_90913,_T_90912,_T_90927,_T_90926,_T_90925,_T_90924,_T_90923,_T_90922}; // @[Mux.scala 19:72:@37407.4]
  assign _T_91750 = {_T_90921,_T_90920,_T_90919,_T_90918,_T_90917,_T_90916,_T_90915,_T_90914,_T_91742}; // @[Mux.scala 19:72:@37415.4]
  assign _T_91752 = _T_90414 ? _T_91750 : 16'h0; // @[Mux.scala 19:72:@37416.4]
  assign _T_91759 = {_T_90984,_T_90999,_T_90998,_T_90997,_T_90996,_T_90995,_T_90994,_T_90993}; // @[Mux.scala 19:72:@37423.4]
  assign _T_91767 = {_T_90992,_T_90991,_T_90990,_T_90989,_T_90988,_T_90987,_T_90986,_T_90985,_T_91759}; // @[Mux.scala 19:72:@37431.4]
  assign _T_91769 = _T_90415 ? _T_91767 : 16'h0; // @[Mux.scala 19:72:@37432.4]
  assign _T_91776 = {_T_91071,_T_91070,_T_91069,_T_91068,_T_91067,_T_91066,_T_91065,_T_91064}; // @[Mux.scala 19:72:@37439.4]
  assign _T_91784 = {_T_91063,_T_91062,_T_91061,_T_91060,_T_91059,_T_91058,_T_91057,_T_91056,_T_91776}; // @[Mux.scala 19:72:@37447.4]
  assign _T_91786 = _T_90416 ? _T_91784 : 16'h0; // @[Mux.scala 19:72:@37448.4]
  assign _T_91793 = {_T_91142,_T_91141,_T_91140,_T_91139,_T_91138,_T_91137,_T_91136,_T_91135}; // @[Mux.scala 19:72:@37455.4]
  assign _T_91801 = {_T_91134,_T_91133,_T_91132,_T_91131,_T_91130,_T_91129,_T_91128,_T_91143,_T_91793}; // @[Mux.scala 19:72:@37463.4]
  assign _T_91803 = _T_90417 ? _T_91801 : 16'h0; // @[Mux.scala 19:72:@37464.4]
  assign _T_91810 = {_T_91213,_T_91212,_T_91211,_T_91210,_T_91209,_T_91208,_T_91207,_T_91206}; // @[Mux.scala 19:72:@37471.4]
  assign _T_91818 = {_T_91205,_T_91204,_T_91203,_T_91202,_T_91201,_T_91200,_T_91215,_T_91214,_T_91810}; // @[Mux.scala 19:72:@37479.4]
  assign _T_91820 = _T_90418 ? _T_91818 : 16'h0; // @[Mux.scala 19:72:@37480.4]
  assign _T_91827 = {_T_91284,_T_91283,_T_91282,_T_91281,_T_91280,_T_91279,_T_91278,_T_91277}; // @[Mux.scala 19:72:@37487.4]
  assign _T_91835 = {_T_91276,_T_91275,_T_91274,_T_91273,_T_91272,_T_91287,_T_91286,_T_91285,_T_91827}; // @[Mux.scala 19:72:@37495.4]
  assign _T_91837 = _T_90419 ? _T_91835 : 16'h0; // @[Mux.scala 19:72:@37496.4]
  assign _T_91844 = {_T_91355,_T_91354,_T_91353,_T_91352,_T_91351,_T_91350,_T_91349,_T_91348}; // @[Mux.scala 19:72:@37503.4]
  assign _T_91852 = {_T_91347,_T_91346,_T_91345,_T_91344,_T_91359,_T_91358,_T_91357,_T_91356,_T_91844}; // @[Mux.scala 19:72:@37511.4]
  assign _T_91854 = _T_90420 ? _T_91852 : 16'h0; // @[Mux.scala 19:72:@37512.4]
  assign _T_91861 = {_T_91426,_T_91425,_T_91424,_T_91423,_T_91422,_T_91421,_T_91420,_T_91419}; // @[Mux.scala 19:72:@37519.4]
  assign _T_91869 = {_T_91418,_T_91417,_T_91416,_T_91431,_T_91430,_T_91429,_T_91428,_T_91427,_T_91861}; // @[Mux.scala 19:72:@37527.4]
  assign _T_91871 = _T_90421 ? _T_91869 : 16'h0; // @[Mux.scala 19:72:@37528.4]
  assign _T_91878 = {_T_91497,_T_91496,_T_91495,_T_91494,_T_91493,_T_91492,_T_91491,_T_91490}; // @[Mux.scala 19:72:@37535.4]
  assign _T_91886 = {_T_91489,_T_91488,_T_91503,_T_91502,_T_91501,_T_91500,_T_91499,_T_91498,_T_91878}; // @[Mux.scala 19:72:@37543.4]
  assign _T_91888 = _T_90422 ? _T_91886 : 16'h0; // @[Mux.scala 19:72:@37544.4]
  assign _T_91895 = {_T_91568,_T_91567,_T_91566,_T_91565,_T_91564,_T_91563,_T_91562,_T_91561}; // @[Mux.scala 19:72:@37551.4]
  assign _T_91903 = {_T_91560,_T_91575,_T_91574,_T_91573,_T_91572,_T_91571,_T_91570,_T_91569,_T_91895}; // @[Mux.scala 19:72:@37559.4]
  assign _T_91905 = _T_90423 ? _T_91903 : 16'h0; // @[Mux.scala 19:72:@37560.4]
  assign _T_91906 = _T_91650 | _T_91667; // @[Mux.scala 19:72:@37561.4]
  assign _T_91907 = _T_91906 | _T_91684; // @[Mux.scala 19:72:@37562.4]
  assign _T_91908 = _T_91907 | _T_91701; // @[Mux.scala 19:72:@37563.4]
  assign _T_91909 = _T_91908 | _T_91718; // @[Mux.scala 19:72:@37564.4]
  assign _T_91910 = _T_91909 | _T_91735; // @[Mux.scala 19:72:@37565.4]
  assign _T_91911 = _T_91910 | _T_91752; // @[Mux.scala 19:72:@37566.4]
  assign _T_91912 = _T_91911 | _T_91769; // @[Mux.scala 19:72:@37567.4]
  assign _T_91913 = _T_91912 | _T_91786; // @[Mux.scala 19:72:@37568.4]
  assign _T_91914 = _T_91913 | _T_91803; // @[Mux.scala 19:72:@37569.4]
  assign _T_91915 = _T_91914 | _T_91820; // @[Mux.scala 19:72:@37570.4]
  assign _T_91916 = _T_91915 | _T_91837; // @[Mux.scala 19:72:@37571.4]
  assign _T_91917 = _T_91916 | _T_91854; // @[Mux.scala 19:72:@37572.4]
  assign _T_91918 = _T_91917 | _T_91871; // @[Mux.scala 19:72:@37573.4]
  assign _T_91919 = _T_91918 | _T_91888; // @[Mux.scala 19:72:@37574.4]
  assign _T_91920 = _T_91919 | _T_91905; // @[Mux.scala 19:72:@37575.4]
  assign priorityLoadRequest_0 = _T_91920[0]; // @[Mux.scala 19:72:@37579.4]
  assign priorityLoadRequest_1 = _T_91920[1]; // @[Mux.scala 19:72:@37581.4]
  assign priorityLoadRequest_2 = _T_91920[2]; // @[Mux.scala 19:72:@37583.4]
  assign priorityLoadRequest_3 = _T_91920[3]; // @[Mux.scala 19:72:@37585.4]
  assign priorityLoadRequest_4 = _T_91920[4]; // @[Mux.scala 19:72:@37587.4]
  assign priorityLoadRequest_5 = _T_91920[5]; // @[Mux.scala 19:72:@37589.4]
  assign priorityLoadRequest_6 = _T_91920[6]; // @[Mux.scala 19:72:@37591.4]
  assign priorityLoadRequest_7 = _T_91920[7]; // @[Mux.scala 19:72:@37593.4]
  assign priorityLoadRequest_8 = _T_91920[8]; // @[Mux.scala 19:72:@37595.4]
  assign priorityLoadRequest_9 = _T_91920[9]; // @[Mux.scala 19:72:@37597.4]
  assign priorityLoadRequest_10 = _T_91920[10]; // @[Mux.scala 19:72:@37599.4]
  assign priorityLoadRequest_11 = _T_91920[11]; // @[Mux.scala 19:72:@37601.4]
  assign priorityLoadRequest_12 = _T_91920[12]; // @[Mux.scala 19:72:@37603.4]
  assign priorityLoadRequest_13 = _T_91920[13]; // @[Mux.scala 19:72:@37605.4]
  assign priorityLoadRequest_14 = _T_91920[14]; // @[Mux.scala 19:72:@37607.4]
  assign priorityLoadRequest_15 = _T_91920[15]; // @[Mux.scala 19:72:@37609.4]
  assign _GEN_1920 = io_memIsReadyForLoads ? priorityLoadRequest_0 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1921 = io_memIsReadyForLoads ? priorityLoadRequest_1 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1922 = io_memIsReadyForLoads ? priorityLoadRequest_2 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1923 = io_memIsReadyForLoads ? priorityLoadRequest_3 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1924 = io_memIsReadyForLoads ? priorityLoadRequest_4 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1925 = io_memIsReadyForLoads ? priorityLoadRequest_5 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1926 = io_memIsReadyForLoads ? priorityLoadRequest_6 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1927 = io_memIsReadyForLoads ? priorityLoadRequest_7 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1928 = io_memIsReadyForLoads ? priorityLoadRequest_8 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1929 = io_memIsReadyForLoads ? priorityLoadRequest_9 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1930 = io_memIsReadyForLoads ? priorityLoadRequest_10 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1931 = io_memIsReadyForLoads ? priorityLoadRequest_11 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1932 = io_memIsReadyForLoads ? priorityLoadRequest_12 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1933 = io_memIsReadyForLoads ? priorityLoadRequest_13 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1934 = io_memIsReadyForLoads ? priorityLoadRequest_14 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1935 = io_memIsReadyForLoads ? priorityLoadRequest_15 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _T_92315 = {storeAddrNotKnownFlagsPReg_0_7,storeAddrNotKnownFlagsPReg_0_6,storeAddrNotKnownFlagsPReg_0_5,storeAddrNotKnownFlagsPReg_0_4,storeAddrNotKnownFlagsPReg_0_3,storeAddrNotKnownFlagsPReg_0_2,storeAddrNotKnownFlagsPReg_0_1,storeAddrNotKnownFlagsPReg_0_0}; // @[LoadQueue.scala 238:58:@37847.8]
  assign _T_92323 = {storeAddrNotKnownFlagsPReg_0_15,storeAddrNotKnownFlagsPReg_0_14,storeAddrNotKnownFlagsPReg_0_13,storeAddrNotKnownFlagsPReg_0_12,storeAddrNotKnownFlagsPReg_0_11,storeAddrNotKnownFlagsPReg_0_10,storeAddrNotKnownFlagsPReg_0_9,storeAddrNotKnownFlagsPReg_0_8,_T_92315}; // @[LoadQueue.scala 238:58:@37855.8]
  assign _T_92330 = {lastConflict_0_7,lastConflict_0_6,lastConflict_0_5,lastConflict_0_4,lastConflict_0_3,lastConflict_0_2,lastConflict_0_1,lastConflict_0_0}; // @[LoadQueue.scala 238:96:@37862.8]
  assign _T_92338 = {lastConflict_0_15,lastConflict_0_14,lastConflict_0_13,lastConflict_0_12,lastConflict_0_11,lastConflict_0_10,lastConflict_0_9,lastConflict_0_8,_T_92330}; // @[LoadQueue.scala 238:96:@37870.8]
  assign _T_92339 = _T_92323 < _T_92338; // @[LoadQueue.scala 238:61:@37871.8]
  assign _T_92340 = canBypass_0 & _T_92339; // @[LoadQueue.scala 237:64:@37872.8]
  assign _GEN_1969 = _T_92269 ? _T_92340 : 1'h0; // @[LoadQueue.scala 230:110:@37804.6]
  assign bypassRequest_0 = _T_92261 ? _GEN_1969 : 1'h0; // @[LoadQueue.scala 229:71:@37798.4]
  assign _GEN_1936 = bypassRequest_0 ? 1'h1 : bypassInitiated_0; // @[LoadQueue.scala 217:34:@37686.6]
  assign _GEN_1937 = initBits_0 ? 1'h0 : _GEN_1936; // @[LoadQueue.scala 215:23:@37682.4]
  assign _T_92399 = {storeAddrNotKnownFlagsPReg_1_7,storeAddrNotKnownFlagsPReg_1_6,storeAddrNotKnownFlagsPReg_1_5,storeAddrNotKnownFlagsPReg_1_4,storeAddrNotKnownFlagsPReg_1_3,storeAddrNotKnownFlagsPReg_1_2,storeAddrNotKnownFlagsPReg_1_1,storeAddrNotKnownFlagsPReg_1_0}; // @[LoadQueue.scala 238:58:@37929.8]
  assign _T_92407 = {storeAddrNotKnownFlagsPReg_1_15,storeAddrNotKnownFlagsPReg_1_14,storeAddrNotKnownFlagsPReg_1_13,storeAddrNotKnownFlagsPReg_1_12,storeAddrNotKnownFlagsPReg_1_11,storeAddrNotKnownFlagsPReg_1_10,storeAddrNotKnownFlagsPReg_1_9,storeAddrNotKnownFlagsPReg_1_8,_T_92399}; // @[LoadQueue.scala 238:58:@37937.8]
  assign _T_92414 = {lastConflict_1_7,lastConflict_1_6,lastConflict_1_5,lastConflict_1_4,lastConflict_1_3,lastConflict_1_2,lastConflict_1_1,lastConflict_1_0}; // @[LoadQueue.scala 238:96:@37944.8]
  assign _T_92422 = {lastConflict_1_15,lastConflict_1_14,lastConflict_1_13,lastConflict_1_12,lastConflict_1_11,lastConflict_1_10,lastConflict_1_9,lastConflict_1_8,_T_92414}; // @[LoadQueue.scala 238:96:@37952.8]
  assign _T_92423 = _T_92407 < _T_92422; // @[LoadQueue.scala 238:61:@37953.8]
  assign _T_92424 = canBypass_1 & _T_92423; // @[LoadQueue.scala 237:64:@37954.8]
  assign _GEN_1973 = _T_92353 ? _T_92424 : 1'h0; // @[LoadQueue.scala 230:110:@37886.6]
  assign bypassRequest_1 = _T_92345 ? _GEN_1973 : 1'h0; // @[LoadQueue.scala 229:71:@37880.4]
  assign _GEN_1938 = bypassRequest_1 ? 1'h1 : bypassInitiated_1; // @[LoadQueue.scala 217:34:@37693.6]
  assign _GEN_1939 = initBits_1 ? 1'h0 : _GEN_1938; // @[LoadQueue.scala 215:23:@37689.4]
  assign _T_92483 = {storeAddrNotKnownFlagsPReg_2_7,storeAddrNotKnownFlagsPReg_2_6,storeAddrNotKnownFlagsPReg_2_5,storeAddrNotKnownFlagsPReg_2_4,storeAddrNotKnownFlagsPReg_2_3,storeAddrNotKnownFlagsPReg_2_2,storeAddrNotKnownFlagsPReg_2_1,storeAddrNotKnownFlagsPReg_2_0}; // @[LoadQueue.scala 238:58:@38011.8]
  assign _T_92491 = {storeAddrNotKnownFlagsPReg_2_15,storeAddrNotKnownFlagsPReg_2_14,storeAddrNotKnownFlagsPReg_2_13,storeAddrNotKnownFlagsPReg_2_12,storeAddrNotKnownFlagsPReg_2_11,storeAddrNotKnownFlagsPReg_2_10,storeAddrNotKnownFlagsPReg_2_9,storeAddrNotKnownFlagsPReg_2_8,_T_92483}; // @[LoadQueue.scala 238:58:@38019.8]
  assign _T_92498 = {lastConflict_2_7,lastConflict_2_6,lastConflict_2_5,lastConflict_2_4,lastConflict_2_3,lastConflict_2_2,lastConflict_2_1,lastConflict_2_0}; // @[LoadQueue.scala 238:96:@38026.8]
  assign _T_92506 = {lastConflict_2_15,lastConflict_2_14,lastConflict_2_13,lastConflict_2_12,lastConflict_2_11,lastConflict_2_10,lastConflict_2_9,lastConflict_2_8,_T_92498}; // @[LoadQueue.scala 238:96:@38034.8]
  assign _T_92507 = _T_92491 < _T_92506; // @[LoadQueue.scala 238:61:@38035.8]
  assign _T_92508 = canBypass_2 & _T_92507; // @[LoadQueue.scala 237:64:@38036.8]
  assign _GEN_1977 = _T_92437 ? _T_92508 : 1'h0; // @[LoadQueue.scala 230:110:@37968.6]
  assign bypassRequest_2 = _T_92429 ? _GEN_1977 : 1'h0; // @[LoadQueue.scala 229:71:@37962.4]
  assign _GEN_1940 = bypassRequest_2 ? 1'h1 : bypassInitiated_2; // @[LoadQueue.scala 217:34:@37700.6]
  assign _GEN_1941 = initBits_2 ? 1'h0 : _GEN_1940; // @[LoadQueue.scala 215:23:@37696.4]
  assign _T_92567 = {storeAddrNotKnownFlagsPReg_3_7,storeAddrNotKnownFlagsPReg_3_6,storeAddrNotKnownFlagsPReg_3_5,storeAddrNotKnownFlagsPReg_3_4,storeAddrNotKnownFlagsPReg_3_3,storeAddrNotKnownFlagsPReg_3_2,storeAddrNotKnownFlagsPReg_3_1,storeAddrNotKnownFlagsPReg_3_0}; // @[LoadQueue.scala 238:58:@38093.8]
  assign _T_92575 = {storeAddrNotKnownFlagsPReg_3_15,storeAddrNotKnownFlagsPReg_3_14,storeAddrNotKnownFlagsPReg_3_13,storeAddrNotKnownFlagsPReg_3_12,storeAddrNotKnownFlagsPReg_3_11,storeAddrNotKnownFlagsPReg_3_10,storeAddrNotKnownFlagsPReg_3_9,storeAddrNotKnownFlagsPReg_3_8,_T_92567}; // @[LoadQueue.scala 238:58:@38101.8]
  assign _T_92582 = {lastConflict_3_7,lastConflict_3_6,lastConflict_3_5,lastConflict_3_4,lastConflict_3_3,lastConflict_3_2,lastConflict_3_1,lastConflict_3_0}; // @[LoadQueue.scala 238:96:@38108.8]
  assign _T_92590 = {lastConflict_3_15,lastConflict_3_14,lastConflict_3_13,lastConflict_3_12,lastConflict_3_11,lastConflict_3_10,lastConflict_3_9,lastConflict_3_8,_T_92582}; // @[LoadQueue.scala 238:96:@38116.8]
  assign _T_92591 = _T_92575 < _T_92590; // @[LoadQueue.scala 238:61:@38117.8]
  assign _T_92592 = canBypass_3 & _T_92591; // @[LoadQueue.scala 237:64:@38118.8]
  assign _GEN_1981 = _T_92521 ? _T_92592 : 1'h0; // @[LoadQueue.scala 230:110:@38050.6]
  assign bypassRequest_3 = _T_92513 ? _GEN_1981 : 1'h0; // @[LoadQueue.scala 229:71:@38044.4]
  assign _GEN_1942 = bypassRequest_3 ? 1'h1 : bypassInitiated_3; // @[LoadQueue.scala 217:34:@37707.6]
  assign _GEN_1943 = initBits_3 ? 1'h0 : _GEN_1942; // @[LoadQueue.scala 215:23:@37703.4]
  assign _T_92651 = {storeAddrNotKnownFlagsPReg_4_7,storeAddrNotKnownFlagsPReg_4_6,storeAddrNotKnownFlagsPReg_4_5,storeAddrNotKnownFlagsPReg_4_4,storeAddrNotKnownFlagsPReg_4_3,storeAddrNotKnownFlagsPReg_4_2,storeAddrNotKnownFlagsPReg_4_1,storeAddrNotKnownFlagsPReg_4_0}; // @[LoadQueue.scala 238:58:@38175.8]
  assign _T_92659 = {storeAddrNotKnownFlagsPReg_4_15,storeAddrNotKnownFlagsPReg_4_14,storeAddrNotKnownFlagsPReg_4_13,storeAddrNotKnownFlagsPReg_4_12,storeAddrNotKnownFlagsPReg_4_11,storeAddrNotKnownFlagsPReg_4_10,storeAddrNotKnownFlagsPReg_4_9,storeAddrNotKnownFlagsPReg_4_8,_T_92651}; // @[LoadQueue.scala 238:58:@38183.8]
  assign _T_92666 = {lastConflict_4_7,lastConflict_4_6,lastConflict_4_5,lastConflict_4_4,lastConflict_4_3,lastConflict_4_2,lastConflict_4_1,lastConflict_4_0}; // @[LoadQueue.scala 238:96:@38190.8]
  assign _T_92674 = {lastConflict_4_15,lastConflict_4_14,lastConflict_4_13,lastConflict_4_12,lastConflict_4_11,lastConflict_4_10,lastConflict_4_9,lastConflict_4_8,_T_92666}; // @[LoadQueue.scala 238:96:@38198.8]
  assign _T_92675 = _T_92659 < _T_92674; // @[LoadQueue.scala 238:61:@38199.8]
  assign _T_92676 = canBypass_4 & _T_92675; // @[LoadQueue.scala 237:64:@38200.8]
  assign _GEN_1985 = _T_92605 ? _T_92676 : 1'h0; // @[LoadQueue.scala 230:110:@38132.6]
  assign bypassRequest_4 = _T_92597 ? _GEN_1985 : 1'h0; // @[LoadQueue.scala 229:71:@38126.4]
  assign _GEN_1944 = bypassRequest_4 ? 1'h1 : bypassInitiated_4; // @[LoadQueue.scala 217:34:@37714.6]
  assign _GEN_1945 = initBits_4 ? 1'h0 : _GEN_1944; // @[LoadQueue.scala 215:23:@37710.4]
  assign _T_92735 = {storeAddrNotKnownFlagsPReg_5_7,storeAddrNotKnownFlagsPReg_5_6,storeAddrNotKnownFlagsPReg_5_5,storeAddrNotKnownFlagsPReg_5_4,storeAddrNotKnownFlagsPReg_5_3,storeAddrNotKnownFlagsPReg_5_2,storeAddrNotKnownFlagsPReg_5_1,storeAddrNotKnownFlagsPReg_5_0}; // @[LoadQueue.scala 238:58:@38257.8]
  assign _T_92743 = {storeAddrNotKnownFlagsPReg_5_15,storeAddrNotKnownFlagsPReg_5_14,storeAddrNotKnownFlagsPReg_5_13,storeAddrNotKnownFlagsPReg_5_12,storeAddrNotKnownFlagsPReg_5_11,storeAddrNotKnownFlagsPReg_5_10,storeAddrNotKnownFlagsPReg_5_9,storeAddrNotKnownFlagsPReg_5_8,_T_92735}; // @[LoadQueue.scala 238:58:@38265.8]
  assign _T_92750 = {lastConflict_5_7,lastConflict_5_6,lastConflict_5_5,lastConflict_5_4,lastConflict_5_3,lastConflict_5_2,lastConflict_5_1,lastConflict_5_0}; // @[LoadQueue.scala 238:96:@38272.8]
  assign _T_92758 = {lastConflict_5_15,lastConflict_5_14,lastConflict_5_13,lastConflict_5_12,lastConflict_5_11,lastConflict_5_10,lastConflict_5_9,lastConflict_5_8,_T_92750}; // @[LoadQueue.scala 238:96:@38280.8]
  assign _T_92759 = _T_92743 < _T_92758; // @[LoadQueue.scala 238:61:@38281.8]
  assign _T_92760 = canBypass_5 & _T_92759; // @[LoadQueue.scala 237:64:@38282.8]
  assign _GEN_1989 = _T_92689 ? _T_92760 : 1'h0; // @[LoadQueue.scala 230:110:@38214.6]
  assign bypassRequest_5 = _T_92681 ? _GEN_1989 : 1'h0; // @[LoadQueue.scala 229:71:@38208.4]
  assign _GEN_1946 = bypassRequest_5 ? 1'h1 : bypassInitiated_5; // @[LoadQueue.scala 217:34:@37721.6]
  assign _GEN_1947 = initBits_5 ? 1'h0 : _GEN_1946; // @[LoadQueue.scala 215:23:@37717.4]
  assign _T_92819 = {storeAddrNotKnownFlagsPReg_6_7,storeAddrNotKnownFlagsPReg_6_6,storeAddrNotKnownFlagsPReg_6_5,storeAddrNotKnownFlagsPReg_6_4,storeAddrNotKnownFlagsPReg_6_3,storeAddrNotKnownFlagsPReg_6_2,storeAddrNotKnownFlagsPReg_6_1,storeAddrNotKnownFlagsPReg_6_0}; // @[LoadQueue.scala 238:58:@38339.8]
  assign _T_92827 = {storeAddrNotKnownFlagsPReg_6_15,storeAddrNotKnownFlagsPReg_6_14,storeAddrNotKnownFlagsPReg_6_13,storeAddrNotKnownFlagsPReg_6_12,storeAddrNotKnownFlagsPReg_6_11,storeAddrNotKnownFlagsPReg_6_10,storeAddrNotKnownFlagsPReg_6_9,storeAddrNotKnownFlagsPReg_6_8,_T_92819}; // @[LoadQueue.scala 238:58:@38347.8]
  assign _T_92834 = {lastConflict_6_7,lastConflict_6_6,lastConflict_6_5,lastConflict_6_4,lastConflict_6_3,lastConflict_6_2,lastConflict_6_1,lastConflict_6_0}; // @[LoadQueue.scala 238:96:@38354.8]
  assign _T_92842 = {lastConflict_6_15,lastConflict_6_14,lastConflict_6_13,lastConflict_6_12,lastConflict_6_11,lastConflict_6_10,lastConflict_6_9,lastConflict_6_8,_T_92834}; // @[LoadQueue.scala 238:96:@38362.8]
  assign _T_92843 = _T_92827 < _T_92842; // @[LoadQueue.scala 238:61:@38363.8]
  assign _T_92844 = canBypass_6 & _T_92843; // @[LoadQueue.scala 237:64:@38364.8]
  assign _GEN_1993 = _T_92773 ? _T_92844 : 1'h0; // @[LoadQueue.scala 230:110:@38296.6]
  assign bypassRequest_6 = _T_92765 ? _GEN_1993 : 1'h0; // @[LoadQueue.scala 229:71:@38290.4]
  assign _GEN_1948 = bypassRequest_6 ? 1'h1 : bypassInitiated_6; // @[LoadQueue.scala 217:34:@37728.6]
  assign _GEN_1949 = initBits_6 ? 1'h0 : _GEN_1948; // @[LoadQueue.scala 215:23:@37724.4]
  assign _T_92903 = {storeAddrNotKnownFlagsPReg_7_7,storeAddrNotKnownFlagsPReg_7_6,storeAddrNotKnownFlagsPReg_7_5,storeAddrNotKnownFlagsPReg_7_4,storeAddrNotKnownFlagsPReg_7_3,storeAddrNotKnownFlagsPReg_7_2,storeAddrNotKnownFlagsPReg_7_1,storeAddrNotKnownFlagsPReg_7_0}; // @[LoadQueue.scala 238:58:@38421.8]
  assign _T_92911 = {storeAddrNotKnownFlagsPReg_7_15,storeAddrNotKnownFlagsPReg_7_14,storeAddrNotKnownFlagsPReg_7_13,storeAddrNotKnownFlagsPReg_7_12,storeAddrNotKnownFlagsPReg_7_11,storeAddrNotKnownFlagsPReg_7_10,storeAddrNotKnownFlagsPReg_7_9,storeAddrNotKnownFlagsPReg_7_8,_T_92903}; // @[LoadQueue.scala 238:58:@38429.8]
  assign _T_92918 = {lastConflict_7_7,lastConflict_7_6,lastConflict_7_5,lastConflict_7_4,lastConflict_7_3,lastConflict_7_2,lastConflict_7_1,lastConflict_7_0}; // @[LoadQueue.scala 238:96:@38436.8]
  assign _T_92926 = {lastConflict_7_15,lastConflict_7_14,lastConflict_7_13,lastConflict_7_12,lastConflict_7_11,lastConflict_7_10,lastConflict_7_9,lastConflict_7_8,_T_92918}; // @[LoadQueue.scala 238:96:@38444.8]
  assign _T_92927 = _T_92911 < _T_92926; // @[LoadQueue.scala 238:61:@38445.8]
  assign _T_92928 = canBypass_7 & _T_92927; // @[LoadQueue.scala 237:64:@38446.8]
  assign _GEN_1997 = _T_92857 ? _T_92928 : 1'h0; // @[LoadQueue.scala 230:110:@38378.6]
  assign bypassRequest_7 = _T_92849 ? _GEN_1997 : 1'h0; // @[LoadQueue.scala 229:71:@38372.4]
  assign _GEN_1950 = bypassRequest_7 ? 1'h1 : bypassInitiated_7; // @[LoadQueue.scala 217:34:@37735.6]
  assign _GEN_1951 = initBits_7 ? 1'h0 : _GEN_1950; // @[LoadQueue.scala 215:23:@37731.4]
  assign _T_92987 = {storeAddrNotKnownFlagsPReg_8_7,storeAddrNotKnownFlagsPReg_8_6,storeAddrNotKnownFlagsPReg_8_5,storeAddrNotKnownFlagsPReg_8_4,storeAddrNotKnownFlagsPReg_8_3,storeAddrNotKnownFlagsPReg_8_2,storeAddrNotKnownFlagsPReg_8_1,storeAddrNotKnownFlagsPReg_8_0}; // @[LoadQueue.scala 238:58:@38503.8]
  assign _T_92995 = {storeAddrNotKnownFlagsPReg_8_15,storeAddrNotKnownFlagsPReg_8_14,storeAddrNotKnownFlagsPReg_8_13,storeAddrNotKnownFlagsPReg_8_12,storeAddrNotKnownFlagsPReg_8_11,storeAddrNotKnownFlagsPReg_8_10,storeAddrNotKnownFlagsPReg_8_9,storeAddrNotKnownFlagsPReg_8_8,_T_92987}; // @[LoadQueue.scala 238:58:@38511.8]
  assign _T_93002 = {lastConflict_8_7,lastConflict_8_6,lastConflict_8_5,lastConflict_8_4,lastConflict_8_3,lastConflict_8_2,lastConflict_8_1,lastConflict_8_0}; // @[LoadQueue.scala 238:96:@38518.8]
  assign _T_93010 = {lastConflict_8_15,lastConflict_8_14,lastConflict_8_13,lastConflict_8_12,lastConflict_8_11,lastConflict_8_10,lastConflict_8_9,lastConflict_8_8,_T_93002}; // @[LoadQueue.scala 238:96:@38526.8]
  assign _T_93011 = _T_92995 < _T_93010; // @[LoadQueue.scala 238:61:@38527.8]
  assign _T_93012 = canBypass_8 & _T_93011; // @[LoadQueue.scala 237:64:@38528.8]
  assign _GEN_2001 = _T_92941 ? _T_93012 : 1'h0; // @[LoadQueue.scala 230:110:@38460.6]
  assign bypassRequest_8 = _T_92933 ? _GEN_2001 : 1'h0; // @[LoadQueue.scala 229:71:@38454.4]
  assign _GEN_1952 = bypassRequest_8 ? 1'h1 : bypassInitiated_8; // @[LoadQueue.scala 217:34:@37742.6]
  assign _GEN_1953 = initBits_8 ? 1'h0 : _GEN_1952; // @[LoadQueue.scala 215:23:@37738.4]
  assign _T_93071 = {storeAddrNotKnownFlagsPReg_9_7,storeAddrNotKnownFlagsPReg_9_6,storeAddrNotKnownFlagsPReg_9_5,storeAddrNotKnownFlagsPReg_9_4,storeAddrNotKnownFlagsPReg_9_3,storeAddrNotKnownFlagsPReg_9_2,storeAddrNotKnownFlagsPReg_9_1,storeAddrNotKnownFlagsPReg_9_0}; // @[LoadQueue.scala 238:58:@38585.8]
  assign _T_93079 = {storeAddrNotKnownFlagsPReg_9_15,storeAddrNotKnownFlagsPReg_9_14,storeAddrNotKnownFlagsPReg_9_13,storeAddrNotKnownFlagsPReg_9_12,storeAddrNotKnownFlagsPReg_9_11,storeAddrNotKnownFlagsPReg_9_10,storeAddrNotKnownFlagsPReg_9_9,storeAddrNotKnownFlagsPReg_9_8,_T_93071}; // @[LoadQueue.scala 238:58:@38593.8]
  assign _T_93086 = {lastConflict_9_7,lastConflict_9_6,lastConflict_9_5,lastConflict_9_4,lastConflict_9_3,lastConflict_9_2,lastConflict_9_1,lastConflict_9_0}; // @[LoadQueue.scala 238:96:@38600.8]
  assign _T_93094 = {lastConflict_9_15,lastConflict_9_14,lastConflict_9_13,lastConflict_9_12,lastConflict_9_11,lastConflict_9_10,lastConflict_9_9,lastConflict_9_8,_T_93086}; // @[LoadQueue.scala 238:96:@38608.8]
  assign _T_93095 = _T_93079 < _T_93094; // @[LoadQueue.scala 238:61:@38609.8]
  assign _T_93096 = canBypass_9 & _T_93095; // @[LoadQueue.scala 237:64:@38610.8]
  assign _GEN_2005 = _T_93025 ? _T_93096 : 1'h0; // @[LoadQueue.scala 230:110:@38542.6]
  assign bypassRequest_9 = _T_93017 ? _GEN_2005 : 1'h0; // @[LoadQueue.scala 229:71:@38536.4]
  assign _GEN_1954 = bypassRequest_9 ? 1'h1 : bypassInitiated_9; // @[LoadQueue.scala 217:34:@37749.6]
  assign _GEN_1955 = initBits_9 ? 1'h0 : _GEN_1954; // @[LoadQueue.scala 215:23:@37745.4]
  assign _T_93155 = {storeAddrNotKnownFlagsPReg_10_7,storeAddrNotKnownFlagsPReg_10_6,storeAddrNotKnownFlagsPReg_10_5,storeAddrNotKnownFlagsPReg_10_4,storeAddrNotKnownFlagsPReg_10_3,storeAddrNotKnownFlagsPReg_10_2,storeAddrNotKnownFlagsPReg_10_1,storeAddrNotKnownFlagsPReg_10_0}; // @[LoadQueue.scala 238:58:@38667.8]
  assign _T_93163 = {storeAddrNotKnownFlagsPReg_10_15,storeAddrNotKnownFlagsPReg_10_14,storeAddrNotKnownFlagsPReg_10_13,storeAddrNotKnownFlagsPReg_10_12,storeAddrNotKnownFlagsPReg_10_11,storeAddrNotKnownFlagsPReg_10_10,storeAddrNotKnownFlagsPReg_10_9,storeAddrNotKnownFlagsPReg_10_8,_T_93155}; // @[LoadQueue.scala 238:58:@38675.8]
  assign _T_93170 = {lastConflict_10_7,lastConflict_10_6,lastConflict_10_5,lastConflict_10_4,lastConflict_10_3,lastConflict_10_2,lastConflict_10_1,lastConflict_10_0}; // @[LoadQueue.scala 238:96:@38682.8]
  assign _T_93178 = {lastConflict_10_15,lastConflict_10_14,lastConflict_10_13,lastConflict_10_12,lastConflict_10_11,lastConflict_10_10,lastConflict_10_9,lastConflict_10_8,_T_93170}; // @[LoadQueue.scala 238:96:@38690.8]
  assign _T_93179 = _T_93163 < _T_93178; // @[LoadQueue.scala 238:61:@38691.8]
  assign _T_93180 = canBypass_10 & _T_93179; // @[LoadQueue.scala 237:64:@38692.8]
  assign _GEN_2009 = _T_93109 ? _T_93180 : 1'h0; // @[LoadQueue.scala 230:110:@38624.6]
  assign bypassRequest_10 = _T_93101 ? _GEN_2009 : 1'h0; // @[LoadQueue.scala 229:71:@38618.4]
  assign _GEN_1956 = bypassRequest_10 ? 1'h1 : bypassInitiated_10; // @[LoadQueue.scala 217:34:@37756.6]
  assign _GEN_1957 = initBits_10 ? 1'h0 : _GEN_1956; // @[LoadQueue.scala 215:23:@37752.4]
  assign _T_93239 = {storeAddrNotKnownFlagsPReg_11_7,storeAddrNotKnownFlagsPReg_11_6,storeAddrNotKnownFlagsPReg_11_5,storeAddrNotKnownFlagsPReg_11_4,storeAddrNotKnownFlagsPReg_11_3,storeAddrNotKnownFlagsPReg_11_2,storeAddrNotKnownFlagsPReg_11_1,storeAddrNotKnownFlagsPReg_11_0}; // @[LoadQueue.scala 238:58:@38749.8]
  assign _T_93247 = {storeAddrNotKnownFlagsPReg_11_15,storeAddrNotKnownFlagsPReg_11_14,storeAddrNotKnownFlagsPReg_11_13,storeAddrNotKnownFlagsPReg_11_12,storeAddrNotKnownFlagsPReg_11_11,storeAddrNotKnownFlagsPReg_11_10,storeAddrNotKnownFlagsPReg_11_9,storeAddrNotKnownFlagsPReg_11_8,_T_93239}; // @[LoadQueue.scala 238:58:@38757.8]
  assign _T_93254 = {lastConflict_11_7,lastConflict_11_6,lastConflict_11_5,lastConflict_11_4,lastConflict_11_3,lastConflict_11_2,lastConflict_11_1,lastConflict_11_0}; // @[LoadQueue.scala 238:96:@38764.8]
  assign _T_93262 = {lastConflict_11_15,lastConflict_11_14,lastConflict_11_13,lastConflict_11_12,lastConflict_11_11,lastConflict_11_10,lastConflict_11_9,lastConflict_11_8,_T_93254}; // @[LoadQueue.scala 238:96:@38772.8]
  assign _T_93263 = _T_93247 < _T_93262; // @[LoadQueue.scala 238:61:@38773.8]
  assign _T_93264 = canBypass_11 & _T_93263; // @[LoadQueue.scala 237:64:@38774.8]
  assign _GEN_2013 = _T_93193 ? _T_93264 : 1'h0; // @[LoadQueue.scala 230:110:@38706.6]
  assign bypassRequest_11 = _T_93185 ? _GEN_2013 : 1'h0; // @[LoadQueue.scala 229:71:@38700.4]
  assign _GEN_1958 = bypassRequest_11 ? 1'h1 : bypassInitiated_11; // @[LoadQueue.scala 217:34:@37763.6]
  assign _GEN_1959 = initBits_11 ? 1'h0 : _GEN_1958; // @[LoadQueue.scala 215:23:@37759.4]
  assign _T_93323 = {storeAddrNotKnownFlagsPReg_12_7,storeAddrNotKnownFlagsPReg_12_6,storeAddrNotKnownFlagsPReg_12_5,storeAddrNotKnownFlagsPReg_12_4,storeAddrNotKnownFlagsPReg_12_3,storeAddrNotKnownFlagsPReg_12_2,storeAddrNotKnownFlagsPReg_12_1,storeAddrNotKnownFlagsPReg_12_0}; // @[LoadQueue.scala 238:58:@38831.8]
  assign _T_93331 = {storeAddrNotKnownFlagsPReg_12_15,storeAddrNotKnownFlagsPReg_12_14,storeAddrNotKnownFlagsPReg_12_13,storeAddrNotKnownFlagsPReg_12_12,storeAddrNotKnownFlagsPReg_12_11,storeAddrNotKnownFlagsPReg_12_10,storeAddrNotKnownFlagsPReg_12_9,storeAddrNotKnownFlagsPReg_12_8,_T_93323}; // @[LoadQueue.scala 238:58:@38839.8]
  assign _T_93338 = {lastConflict_12_7,lastConflict_12_6,lastConflict_12_5,lastConflict_12_4,lastConflict_12_3,lastConflict_12_2,lastConflict_12_1,lastConflict_12_0}; // @[LoadQueue.scala 238:96:@38846.8]
  assign _T_93346 = {lastConflict_12_15,lastConflict_12_14,lastConflict_12_13,lastConflict_12_12,lastConflict_12_11,lastConflict_12_10,lastConflict_12_9,lastConflict_12_8,_T_93338}; // @[LoadQueue.scala 238:96:@38854.8]
  assign _T_93347 = _T_93331 < _T_93346; // @[LoadQueue.scala 238:61:@38855.8]
  assign _T_93348 = canBypass_12 & _T_93347; // @[LoadQueue.scala 237:64:@38856.8]
  assign _GEN_2017 = _T_93277 ? _T_93348 : 1'h0; // @[LoadQueue.scala 230:110:@38788.6]
  assign bypassRequest_12 = _T_93269 ? _GEN_2017 : 1'h0; // @[LoadQueue.scala 229:71:@38782.4]
  assign _GEN_1960 = bypassRequest_12 ? 1'h1 : bypassInitiated_12; // @[LoadQueue.scala 217:34:@37770.6]
  assign _GEN_1961 = initBits_12 ? 1'h0 : _GEN_1960; // @[LoadQueue.scala 215:23:@37766.4]
  assign _T_93407 = {storeAddrNotKnownFlagsPReg_13_7,storeAddrNotKnownFlagsPReg_13_6,storeAddrNotKnownFlagsPReg_13_5,storeAddrNotKnownFlagsPReg_13_4,storeAddrNotKnownFlagsPReg_13_3,storeAddrNotKnownFlagsPReg_13_2,storeAddrNotKnownFlagsPReg_13_1,storeAddrNotKnownFlagsPReg_13_0}; // @[LoadQueue.scala 238:58:@38913.8]
  assign _T_93415 = {storeAddrNotKnownFlagsPReg_13_15,storeAddrNotKnownFlagsPReg_13_14,storeAddrNotKnownFlagsPReg_13_13,storeAddrNotKnownFlagsPReg_13_12,storeAddrNotKnownFlagsPReg_13_11,storeAddrNotKnownFlagsPReg_13_10,storeAddrNotKnownFlagsPReg_13_9,storeAddrNotKnownFlagsPReg_13_8,_T_93407}; // @[LoadQueue.scala 238:58:@38921.8]
  assign _T_93422 = {lastConflict_13_7,lastConflict_13_6,lastConflict_13_5,lastConflict_13_4,lastConflict_13_3,lastConflict_13_2,lastConflict_13_1,lastConflict_13_0}; // @[LoadQueue.scala 238:96:@38928.8]
  assign _T_93430 = {lastConflict_13_15,lastConflict_13_14,lastConflict_13_13,lastConflict_13_12,lastConflict_13_11,lastConflict_13_10,lastConflict_13_9,lastConflict_13_8,_T_93422}; // @[LoadQueue.scala 238:96:@38936.8]
  assign _T_93431 = _T_93415 < _T_93430; // @[LoadQueue.scala 238:61:@38937.8]
  assign _T_93432 = canBypass_13 & _T_93431; // @[LoadQueue.scala 237:64:@38938.8]
  assign _GEN_2021 = _T_93361 ? _T_93432 : 1'h0; // @[LoadQueue.scala 230:110:@38870.6]
  assign bypassRequest_13 = _T_93353 ? _GEN_2021 : 1'h0; // @[LoadQueue.scala 229:71:@38864.4]
  assign _GEN_1962 = bypassRequest_13 ? 1'h1 : bypassInitiated_13; // @[LoadQueue.scala 217:34:@37777.6]
  assign _GEN_1963 = initBits_13 ? 1'h0 : _GEN_1962; // @[LoadQueue.scala 215:23:@37773.4]
  assign _T_93491 = {storeAddrNotKnownFlagsPReg_14_7,storeAddrNotKnownFlagsPReg_14_6,storeAddrNotKnownFlagsPReg_14_5,storeAddrNotKnownFlagsPReg_14_4,storeAddrNotKnownFlagsPReg_14_3,storeAddrNotKnownFlagsPReg_14_2,storeAddrNotKnownFlagsPReg_14_1,storeAddrNotKnownFlagsPReg_14_0}; // @[LoadQueue.scala 238:58:@38995.8]
  assign _T_93499 = {storeAddrNotKnownFlagsPReg_14_15,storeAddrNotKnownFlagsPReg_14_14,storeAddrNotKnownFlagsPReg_14_13,storeAddrNotKnownFlagsPReg_14_12,storeAddrNotKnownFlagsPReg_14_11,storeAddrNotKnownFlagsPReg_14_10,storeAddrNotKnownFlagsPReg_14_9,storeAddrNotKnownFlagsPReg_14_8,_T_93491}; // @[LoadQueue.scala 238:58:@39003.8]
  assign _T_93506 = {lastConflict_14_7,lastConflict_14_6,lastConflict_14_5,lastConflict_14_4,lastConflict_14_3,lastConflict_14_2,lastConflict_14_1,lastConflict_14_0}; // @[LoadQueue.scala 238:96:@39010.8]
  assign _T_93514 = {lastConflict_14_15,lastConflict_14_14,lastConflict_14_13,lastConflict_14_12,lastConflict_14_11,lastConflict_14_10,lastConflict_14_9,lastConflict_14_8,_T_93506}; // @[LoadQueue.scala 238:96:@39018.8]
  assign _T_93515 = _T_93499 < _T_93514; // @[LoadQueue.scala 238:61:@39019.8]
  assign _T_93516 = canBypass_14 & _T_93515; // @[LoadQueue.scala 237:64:@39020.8]
  assign _GEN_2025 = _T_93445 ? _T_93516 : 1'h0; // @[LoadQueue.scala 230:110:@38952.6]
  assign bypassRequest_14 = _T_93437 ? _GEN_2025 : 1'h0; // @[LoadQueue.scala 229:71:@38946.4]
  assign _GEN_1964 = bypassRequest_14 ? 1'h1 : bypassInitiated_14; // @[LoadQueue.scala 217:34:@37784.6]
  assign _GEN_1965 = initBits_14 ? 1'h0 : _GEN_1964; // @[LoadQueue.scala 215:23:@37780.4]
  assign _T_93575 = {storeAddrNotKnownFlagsPReg_15_7,storeAddrNotKnownFlagsPReg_15_6,storeAddrNotKnownFlagsPReg_15_5,storeAddrNotKnownFlagsPReg_15_4,storeAddrNotKnownFlagsPReg_15_3,storeAddrNotKnownFlagsPReg_15_2,storeAddrNotKnownFlagsPReg_15_1,storeAddrNotKnownFlagsPReg_15_0}; // @[LoadQueue.scala 238:58:@39077.8]
  assign _T_93583 = {storeAddrNotKnownFlagsPReg_15_15,storeAddrNotKnownFlagsPReg_15_14,storeAddrNotKnownFlagsPReg_15_13,storeAddrNotKnownFlagsPReg_15_12,storeAddrNotKnownFlagsPReg_15_11,storeAddrNotKnownFlagsPReg_15_10,storeAddrNotKnownFlagsPReg_15_9,storeAddrNotKnownFlagsPReg_15_8,_T_93575}; // @[LoadQueue.scala 238:58:@39085.8]
  assign _T_93590 = {lastConflict_15_7,lastConflict_15_6,lastConflict_15_5,lastConflict_15_4,lastConflict_15_3,lastConflict_15_2,lastConflict_15_1,lastConflict_15_0}; // @[LoadQueue.scala 238:96:@39092.8]
  assign _T_93598 = {lastConflict_15_15,lastConflict_15_14,lastConflict_15_13,lastConflict_15_12,lastConflict_15_11,lastConflict_15_10,lastConflict_15_9,lastConflict_15_8,_T_93590}; // @[LoadQueue.scala 238:96:@39100.8]
  assign _T_93599 = _T_93583 < _T_93598; // @[LoadQueue.scala 238:61:@39101.8]
  assign _T_93600 = canBypass_15 & _T_93599; // @[LoadQueue.scala 237:64:@39102.8]
  assign _GEN_2029 = _T_93529 ? _T_93600 : 1'h0; // @[LoadQueue.scala 230:110:@39034.6]
  assign bypassRequest_15 = _T_93521 ? _GEN_2029 : 1'h0; // @[LoadQueue.scala 229:71:@39028.4]
  assign _GEN_1966 = bypassRequest_15 ? 1'h1 : bypassInitiated_15; // @[LoadQueue.scala 217:34:@37791.6]
  assign _GEN_1967 = initBits_15 ? 1'h0 : _GEN_1966; // @[LoadQueue.scala 215:23:@37787.4]
  assign _T_93604 = loadRequest_0 | loadRequest_1; // @[LoadQueue.scala 247:28:@39108.4]
  assign _T_93605 = _T_93604 | loadRequest_2; // @[LoadQueue.scala 247:28:@39109.4]
  assign _T_93606 = _T_93605 | loadRequest_3; // @[LoadQueue.scala 247:28:@39110.4]
  assign _T_93607 = _T_93606 | loadRequest_4; // @[LoadQueue.scala 247:28:@39111.4]
  assign _T_93608 = _T_93607 | loadRequest_5; // @[LoadQueue.scala 247:28:@39112.4]
  assign _T_93609 = _T_93608 | loadRequest_6; // @[LoadQueue.scala 247:28:@39113.4]
  assign _T_93610 = _T_93609 | loadRequest_7; // @[LoadQueue.scala 247:28:@39114.4]
  assign _T_93611 = _T_93610 | loadRequest_8; // @[LoadQueue.scala 247:28:@39115.4]
  assign _T_93612 = _T_93611 | loadRequest_9; // @[LoadQueue.scala 247:28:@39116.4]
  assign _T_93613 = _T_93612 | loadRequest_10; // @[LoadQueue.scala 247:28:@39117.4]
  assign _T_93614 = _T_93613 | loadRequest_11; // @[LoadQueue.scala 247:28:@39118.4]
  assign _T_93615 = _T_93614 | loadRequest_12; // @[LoadQueue.scala 247:28:@39119.4]
  assign _T_93616 = _T_93615 | loadRequest_13; // @[LoadQueue.scala 247:28:@39120.4]
  assign _T_93617 = _T_93616 | loadRequest_14; // @[LoadQueue.scala 247:28:@39121.4]
  assign _T_93618 = _T_93617 | loadRequest_15; // @[LoadQueue.scala 247:28:@39122.4]
  assign _T_93635 = priorityLoadRequest_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@39124.6]
  assign _T_93636 = priorityLoadRequest_13 ? 4'hd : _T_93635; // @[Mux.scala 31:69:@39125.6]
  assign _T_93637 = priorityLoadRequest_12 ? 4'hc : _T_93636; // @[Mux.scala 31:69:@39126.6]
  assign _T_93638 = priorityLoadRequest_11 ? 4'hb : _T_93637; // @[Mux.scala 31:69:@39127.6]
  assign _T_93639 = priorityLoadRequest_10 ? 4'ha : _T_93638; // @[Mux.scala 31:69:@39128.6]
  assign _T_93640 = priorityLoadRequest_9 ? 4'h9 : _T_93639; // @[Mux.scala 31:69:@39129.6]
  assign _T_93641 = priorityLoadRequest_8 ? 4'h8 : _T_93640; // @[Mux.scala 31:69:@39130.6]
  assign _T_93642 = priorityLoadRequest_7 ? 4'h7 : _T_93641; // @[Mux.scala 31:69:@39131.6]
  assign _T_93643 = priorityLoadRequest_6 ? 4'h6 : _T_93642; // @[Mux.scala 31:69:@39132.6]
  assign _T_93644 = priorityLoadRequest_5 ? 4'h5 : _T_93643; // @[Mux.scala 31:69:@39133.6]
  assign _T_93645 = priorityLoadRequest_4 ? 4'h4 : _T_93644; // @[Mux.scala 31:69:@39134.6]
  assign _T_93646 = priorityLoadRequest_3 ? 4'h3 : _T_93645; // @[Mux.scala 31:69:@39135.6]
  assign _T_93647 = priorityLoadRequest_2 ? 4'h2 : _T_93646; // @[Mux.scala 31:69:@39136.6]
  assign _T_93648 = priorityLoadRequest_1 ? 4'h1 : _T_93647; // @[Mux.scala 31:69:@39137.6]
  assign _T_93649 = priorityLoadRequest_0 ? 4'h0 : _T_93648; // @[Mux.scala 31:69:@39138.6]
  assign _GEN_2033 = 4'h1 == _T_93649 ? addrQ_1 : addrQ_0; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2034 = 4'h2 == _T_93649 ? addrQ_2 : _GEN_2033; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2035 = 4'h3 == _T_93649 ? addrQ_3 : _GEN_2034; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2036 = 4'h4 == _T_93649 ? addrQ_4 : _GEN_2035; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2037 = 4'h5 == _T_93649 ? addrQ_5 : _GEN_2036; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2038 = 4'h6 == _T_93649 ? addrQ_6 : _GEN_2037; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2039 = 4'h7 == _T_93649 ? addrQ_7 : _GEN_2038; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2040 = 4'h8 == _T_93649 ? addrQ_8 : _GEN_2039; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2041 = 4'h9 == _T_93649 ? addrQ_9 : _GEN_2040; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2042 = 4'ha == _T_93649 ? addrQ_10 : _GEN_2041; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2043 = 4'hb == _T_93649 ? addrQ_11 : _GEN_2042; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2044 = 4'hc == _T_93649 ? addrQ_12 : _GEN_2043; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2045 = 4'hd == _T_93649 ? addrQ_13 : _GEN_2044; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2046 = 4'he == _T_93649 ? addrQ_14 : _GEN_2045; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2047 = 4'hf == _T_93649 ? addrQ_15 : _GEN_2046; // @[LoadQueue.scala 248:24:@39139.6]
  assign _T_93657 = prevPriorityRequest_0 | bypassRequest_0; // @[LoadQueue.scala 261:41:@39150.6]
  assign _GEN_2050 = _T_93657 ? 1'h1 : dataKnown_0; // @[LoadQueue.scala 261:62:@39151.6]
  assign _GEN_2051 = initBits_0 ? 1'h0 : _GEN_2050; // @[LoadQueue.scala 259:25:@39146.4]
  assign _T_93660 = prevPriorityRequest_1 | bypassRequest_1; // @[LoadQueue.scala 261:41:@39158.6]
  assign _GEN_2052 = _T_93660 ? 1'h1 : dataKnown_1; // @[LoadQueue.scala 261:62:@39159.6]
  assign _GEN_2053 = initBits_1 ? 1'h0 : _GEN_2052; // @[LoadQueue.scala 259:25:@39154.4]
  assign _T_93663 = prevPriorityRequest_2 | bypassRequest_2; // @[LoadQueue.scala 261:41:@39166.6]
  assign _GEN_2054 = _T_93663 ? 1'h1 : dataKnown_2; // @[LoadQueue.scala 261:62:@39167.6]
  assign _GEN_2055 = initBits_2 ? 1'h0 : _GEN_2054; // @[LoadQueue.scala 259:25:@39162.4]
  assign _T_93666 = prevPriorityRequest_3 | bypassRequest_3; // @[LoadQueue.scala 261:41:@39174.6]
  assign _GEN_2056 = _T_93666 ? 1'h1 : dataKnown_3; // @[LoadQueue.scala 261:62:@39175.6]
  assign _GEN_2057 = initBits_3 ? 1'h0 : _GEN_2056; // @[LoadQueue.scala 259:25:@39170.4]
  assign _T_93669 = prevPriorityRequest_4 | bypassRequest_4; // @[LoadQueue.scala 261:41:@39182.6]
  assign _GEN_2058 = _T_93669 ? 1'h1 : dataKnown_4; // @[LoadQueue.scala 261:62:@39183.6]
  assign _GEN_2059 = initBits_4 ? 1'h0 : _GEN_2058; // @[LoadQueue.scala 259:25:@39178.4]
  assign _T_93672 = prevPriorityRequest_5 | bypassRequest_5; // @[LoadQueue.scala 261:41:@39190.6]
  assign _GEN_2060 = _T_93672 ? 1'h1 : dataKnown_5; // @[LoadQueue.scala 261:62:@39191.6]
  assign _GEN_2061 = initBits_5 ? 1'h0 : _GEN_2060; // @[LoadQueue.scala 259:25:@39186.4]
  assign _T_93675 = prevPriorityRequest_6 | bypassRequest_6; // @[LoadQueue.scala 261:41:@39198.6]
  assign _GEN_2062 = _T_93675 ? 1'h1 : dataKnown_6; // @[LoadQueue.scala 261:62:@39199.6]
  assign _GEN_2063 = initBits_6 ? 1'h0 : _GEN_2062; // @[LoadQueue.scala 259:25:@39194.4]
  assign _T_93678 = prevPriorityRequest_7 | bypassRequest_7; // @[LoadQueue.scala 261:41:@39206.6]
  assign _GEN_2064 = _T_93678 ? 1'h1 : dataKnown_7; // @[LoadQueue.scala 261:62:@39207.6]
  assign _GEN_2065 = initBits_7 ? 1'h0 : _GEN_2064; // @[LoadQueue.scala 259:25:@39202.4]
  assign _T_93681 = prevPriorityRequest_8 | bypassRequest_8; // @[LoadQueue.scala 261:41:@39214.6]
  assign _GEN_2066 = _T_93681 ? 1'h1 : dataKnown_8; // @[LoadQueue.scala 261:62:@39215.6]
  assign _GEN_2067 = initBits_8 ? 1'h0 : _GEN_2066; // @[LoadQueue.scala 259:25:@39210.4]
  assign _T_93684 = prevPriorityRequest_9 | bypassRequest_9; // @[LoadQueue.scala 261:41:@39222.6]
  assign _GEN_2068 = _T_93684 ? 1'h1 : dataKnown_9; // @[LoadQueue.scala 261:62:@39223.6]
  assign _GEN_2069 = initBits_9 ? 1'h0 : _GEN_2068; // @[LoadQueue.scala 259:25:@39218.4]
  assign _T_93687 = prevPriorityRequest_10 | bypassRequest_10; // @[LoadQueue.scala 261:41:@39230.6]
  assign _GEN_2070 = _T_93687 ? 1'h1 : dataKnown_10; // @[LoadQueue.scala 261:62:@39231.6]
  assign _GEN_2071 = initBits_10 ? 1'h0 : _GEN_2070; // @[LoadQueue.scala 259:25:@39226.4]
  assign _T_93690 = prevPriorityRequest_11 | bypassRequest_11; // @[LoadQueue.scala 261:41:@39238.6]
  assign _GEN_2072 = _T_93690 ? 1'h1 : dataKnown_11; // @[LoadQueue.scala 261:62:@39239.6]
  assign _GEN_2073 = initBits_11 ? 1'h0 : _GEN_2072; // @[LoadQueue.scala 259:25:@39234.4]
  assign _T_93693 = prevPriorityRequest_12 | bypassRequest_12; // @[LoadQueue.scala 261:41:@39246.6]
  assign _GEN_2074 = _T_93693 ? 1'h1 : dataKnown_12; // @[LoadQueue.scala 261:62:@39247.6]
  assign _GEN_2075 = initBits_12 ? 1'h0 : _GEN_2074; // @[LoadQueue.scala 259:25:@39242.4]
  assign _T_93696 = prevPriorityRequest_13 | bypassRequest_13; // @[LoadQueue.scala 261:41:@39254.6]
  assign _GEN_2076 = _T_93696 ? 1'h1 : dataKnown_13; // @[LoadQueue.scala 261:62:@39255.6]
  assign _GEN_2077 = initBits_13 ? 1'h0 : _GEN_2076; // @[LoadQueue.scala 259:25:@39250.4]
  assign _T_93699 = prevPriorityRequest_14 | bypassRequest_14; // @[LoadQueue.scala 261:41:@39262.6]
  assign _GEN_2078 = _T_93699 ? 1'h1 : dataKnown_14; // @[LoadQueue.scala 261:62:@39263.6]
  assign _GEN_2079 = initBits_14 ? 1'h0 : _GEN_2078; // @[LoadQueue.scala 259:25:@39258.4]
  assign _T_93702 = prevPriorityRequest_15 | bypassRequest_15; // @[LoadQueue.scala 261:41:@39270.6]
  assign _GEN_2080 = _T_93702 ? 1'h1 : dataKnown_15; // @[LoadQueue.scala 261:62:@39271.6]
  assign _GEN_2081 = initBits_15 ? 1'h0 : _GEN_2080; // @[LoadQueue.scala 259:25:@39266.4]
  assign _GEN_2082 = prevPriorityRequest_0 ? io_loadDataFromMem : dataQ_0; // @[LoadQueue.scala 269:44:@39278.6]
  assign _GEN_2083 = bypassRequest_0 ? bypassVal_0 : _GEN_2082; // @[LoadQueue.scala 267:32:@39274.4]
  assign _GEN_2084 = prevPriorityRequest_1 ? io_loadDataFromMem : dataQ_1; // @[LoadQueue.scala 269:44:@39285.6]
  assign _GEN_2085 = bypassRequest_1 ? bypassVal_1 : _GEN_2084; // @[LoadQueue.scala 267:32:@39281.4]
  assign _GEN_2086 = prevPriorityRequest_2 ? io_loadDataFromMem : dataQ_2; // @[LoadQueue.scala 269:44:@39292.6]
  assign _GEN_2087 = bypassRequest_2 ? bypassVal_2 : _GEN_2086; // @[LoadQueue.scala 267:32:@39288.4]
  assign _GEN_2088 = prevPriorityRequest_3 ? io_loadDataFromMem : dataQ_3; // @[LoadQueue.scala 269:44:@39299.6]
  assign _GEN_2089 = bypassRequest_3 ? bypassVal_3 : _GEN_2088; // @[LoadQueue.scala 267:32:@39295.4]
  assign _GEN_2090 = prevPriorityRequest_4 ? io_loadDataFromMem : dataQ_4; // @[LoadQueue.scala 269:44:@39306.6]
  assign _GEN_2091 = bypassRequest_4 ? bypassVal_4 : _GEN_2090; // @[LoadQueue.scala 267:32:@39302.4]
  assign _GEN_2092 = prevPriorityRequest_5 ? io_loadDataFromMem : dataQ_5; // @[LoadQueue.scala 269:44:@39313.6]
  assign _GEN_2093 = bypassRequest_5 ? bypassVal_5 : _GEN_2092; // @[LoadQueue.scala 267:32:@39309.4]
  assign _GEN_2094 = prevPriorityRequest_6 ? io_loadDataFromMem : dataQ_6; // @[LoadQueue.scala 269:44:@39320.6]
  assign _GEN_2095 = bypassRequest_6 ? bypassVal_6 : _GEN_2094; // @[LoadQueue.scala 267:32:@39316.4]
  assign _GEN_2096 = prevPriorityRequest_7 ? io_loadDataFromMem : dataQ_7; // @[LoadQueue.scala 269:44:@39327.6]
  assign _GEN_2097 = bypassRequest_7 ? bypassVal_7 : _GEN_2096; // @[LoadQueue.scala 267:32:@39323.4]
  assign _GEN_2098 = prevPriorityRequest_8 ? io_loadDataFromMem : dataQ_8; // @[LoadQueue.scala 269:44:@39334.6]
  assign _GEN_2099 = bypassRequest_8 ? bypassVal_8 : _GEN_2098; // @[LoadQueue.scala 267:32:@39330.4]
  assign _GEN_2100 = prevPriorityRequest_9 ? io_loadDataFromMem : dataQ_9; // @[LoadQueue.scala 269:44:@39341.6]
  assign _GEN_2101 = bypassRequest_9 ? bypassVal_9 : _GEN_2100; // @[LoadQueue.scala 267:32:@39337.4]
  assign _GEN_2102 = prevPriorityRequest_10 ? io_loadDataFromMem : dataQ_10; // @[LoadQueue.scala 269:44:@39348.6]
  assign _GEN_2103 = bypassRequest_10 ? bypassVal_10 : _GEN_2102; // @[LoadQueue.scala 267:32:@39344.4]
  assign _GEN_2104 = prevPriorityRequest_11 ? io_loadDataFromMem : dataQ_11; // @[LoadQueue.scala 269:44:@39355.6]
  assign _GEN_2105 = bypassRequest_11 ? bypassVal_11 : _GEN_2104; // @[LoadQueue.scala 267:32:@39351.4]
  assign _GEN_2106 = prevPriorityRequest_12 ? io_loadDataFromMem : dataQ_12; // @[LoadQueue.scala 269:44:@39362.6]
  assign _GEN_2107 = bypassRequest_12 ? bypassVal_12 : _GEN_2106; // @[LoadQueue.scala 267:32:@39358.4]
  assign _GEN_2108 = prevPriorityRequest_13 ? io_loadDataFromMem : dataQ_13; // @[LoadQueue.scala 269:44:@39369.6]
  assign _GEN_2109 = bypassRequest_13 ? bypassVal_13 : _GEN_2108; // @[LoadQueue.scala 267:32:@39365.4]
  assign _GEN_2110 = prevPriorityRequest_14 ? io_loadDataFromMem : dataQ_14; // @[LoadQueue.scala 269:44:@39376.6]
  assign _GEN_2111 = bypassRequest_14 ? bypassVal_14 : _GEN_2110; // @[LoadQueue.scala 267:32:@39372.4]
  assign _GEN_2112 = prevPriorityRequest_15 ? io_loadDataFromMem : dataQ_15; // @[LoadQueue.scala 269:44:@39383.6]
  assign _GEN_2113 = bypassRequest_15 ? bypassVal_15 : _GEN_2112; // @[LoadQueue.scala 267:32:@39379.4]
  assign entriesPorts_0_0 = portQ_0 == 1'h0; // @[LoadQueue.scala 286:69:@39387.4]
  assign entriesPorts_0_1 = portQ_1 == 1'h0; // @[LoadQueue.scala 286:69:@39389.4]
  assign entriesPorts_0_2 = portQ_2 == 1'h0; // @[LoadQueue.scala 286:69:@39391.4]
  assign entriesPorts_0_3 = portQ_3 == 1'h0; // @[LoadQueue.scala 286:69:@39393.4]
  assign entriesPorts_0_4 = portQ_4 == 1'h0; // @[LoadQueue.scala 286:69:@39395.4]
  assign entriesPorts_0_5 = portQ_5 == 1'h0; // @[LoadQueue.scala 286:69:@39397.4]
  assign entriesPorts_0_6 = portQ_6 == 1'h0; // @[LoadQueue.scala 286:69:@39399.4]
  assign entriesPorts_0_7 = portQ_7 == 1'h0; // @[LoadQueue.scala 286:69:@39401.4]
  assign entriesPorts_0_8 = portQ_8 == 1'h0; // @[LoadQueue.scala 286:69:@39403.4]
  assign entriesPorts_0_9 = portQ_9 == 1'h0; // @[LoadQueue.scala 286:69:@39405.4]
  assign entriesPorts_0_10 = portQ_10 == 1'h0; // @[LoadQueue.scala 286:69:@39407.4]
  assign entriesPorts_0_11 = portQ_11 == 1'h0; // @[LoadQueue.scala 286:69:@39409.4]
  assign entriesPorts_0_12 = portQ_12 == 1'h0; // @[LoadQueue.scala 286:69:@39411.4]
  assign entriesPorts_0_13 = portQ_13 == 1'h0; // @[LoadQueue.scala 286:69:@39413.4]
  assign entriesPorts_0_14 = portQ_14 == 1'h0; // @[LoadQueue.scala 286:69:@39415.4]
  assign entriesPorts_0_15 = portQ_15 == 1'h0; // @[LoadQueue.scala 286:69:@39417.4]
  assign _T_94435 = addrKnown_0 == 1'h0; // @[LoadQueue.scala 298:86:@39453.4]
  assign _T_94436 = entriesPorts_0_0 & _T_94435; // @[LoadQueue.scala 298:83:@39454.4]
  assign _T_94438 = addrKnown_1 == 1'h0; // @[LoadQueue.scala 298:86:@39455.4]
  assign _T_94439 = entriesPorts_0_1 & _T_94438; // @[LoadQueue.scala 298:83:@39456.4]
  assign _T_94441 = addrKnown_2 == 1'h0; // @[LoadQueue.scala 298:86:@39457.4]
  assign _T_94442 = entriesPorts_0_2 & _T_94441; // @[LoadQueue.scala 298:83:@39458.4]
  assign _T_94444 = addrKnown_3 == 1'h0; // @[LoadQueue.scala 298:86:@39459.4]
  assign _T_94445 = entriesPorts_0_3 & _T_94444; // @[LoadQueue.scala 298:83:@39460.4]
  assign _T_94447 = addrKnown_4 == 1'h0; // @[LoadQueue.scala 298:86:@39461.4]
  assign _T_94448 = entriesPorts_0_4 & _T_94447; // @[LoadQueue.scala 298:83:@39462.4]
  assign _T_94450 = addrKnown_5 == 1'h0; // @[LoadQueue.scala 298:86:@39463.4]
  assign _T_94451 = entriesPorts_0_5 & _T_94450; // @[LoadQueue.scala 298:83:@39464.4]
  assign _T_94453 = addrKnown_6 == 1'h0; // @[LoadQueue.scala 298:86:@39465.4]
  assign _T_94454 = entriesPorts_0_6 & _T_94453; // @[LoadQueue.scala 298:83:@39466.4]
  assign _T_94456 = addrKnown_7 == 1'h0; // @[LoadQueue.scala 298:86:@39467.4]
  assign _T_94457 = entriesPorts_0_7 & _T_94456; // @[LoadQueue.scala 298:83:@39468.4]
  assign _T_94459 = addrKnown_8 == 1'h0; // @[LoadQueue.scala 298:86:@39469.4]
  assign _T_94460 = entriesPorts_0_8 & _T_94459; // @[LoadQueue.scala 298:83:@39470.4]
  assign _T_94462 = addrKnown_9 == 1'h0; // @[LoadQueue.scala 298:86:@39471.4]
  assign _T_94463 = entriesPorts_0_9 & _T_94462; // @[LoadQueue.scala 298:83:@39472.4]
  assign _T_94465 = addrKnown_10 == 1'h0; // @[LoadQueue.scala 298:86:@39473.4]
  assign _T_94466 = entriesPorts_0_10 & _T_94465; // @[LoadQueue.scala 298:83:@39474.4]
  assign _T_94468 = addrKnown_11 == 1'h0; // @[LoadQueue.scala 298:86:@39475.4]
  assign _T_94469 = entriesPorts_0_11 & _T_94468; // @[LoadQueue.scala 298:83:@39476.4]
  assign _T_94471 = addrKnown_12 == 1'h0; // @[LoadQueue.scala 298:86:@39477.4]
  assign _T_94472 = entriesPorts_0_12 & _T_94471; // @[LoadQueue.scala 298:83:@39478.4]
  assign _T_94474 = addrKnown_13 == 1'h0; // @[LoadQueue.scala 298:86:@39479.4]
  assign _T_94475 = entriesPorts_0_13 & _T_94474; // @[LoadQueue.scala 298:83:@39480.4]
  assign _T_94477 = addrKnown_14 == 1'h0; // @[LoadQueue.scala 298:86:@39481.4]
  assign _T_94478 = entriesPorts_0_14 & _T_94477; // @[LoadQueue.scala 298:83:@39482.4]
  assign _T_94480 = addrKnown_15 == 1'h0; // @[LoadQueue.scala 298:86:@39483.4]
  assign _T_94481 = entriesPorts_0_15 & _T_94480; // @[LoadQueue.scala 298:83:@39484.4]
  assign _T_94564 = _T_94481 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39538.4]
  assign _T_94565 = _T_94478 ? 16'h4000 : _T_94564; // @[Mux.scala 31:69:@39539.4]
  assign _T_94566 = _T_94475 ? 16'h2000 : _T_94565; // @[Mux.scala 31:69:@39540.4]
  assign _T_94567 = _T_94472 ? 16'h1000 : _T_94566; // @[Mux.scala 31:69:@39541.4]
  assign _T_94568 = _T_94469 ? 16'h800 : _T_94567; // @[Mux.scala 31:69:@39542.4]
  assign _T_94569 = _T_94466 ? 16'h400 : _T_94568; // @[Mux.scala 31:69:@39543.4]
  assign _T_94570 = _T_94463 ? 16'h200 : _T_94569; // @[Mux.scala 31:69:@39544.4]
  assign _T_94571 = _T_94460 ? 16'h100 : _T_94570; // @[Mux.scala 31:69:@39545.4]
  assign _T_94572 = _T_94457 ? 16'h80 : _T_94571; // @[Mux.scala 31:69:@39546.4]
  assign _T_94573 = _T_94454 ? 16'h40 : _T_94572; // @[Mux.scala 31:69:@39547.4]
  assign _T_94574 = _T_94451 ? 16'h20 : _T_94573; // @[Mux.scala 31:69:@39548.4]
  assign _T_94575 = _T_94448 ? 16'h10 : _T_94574; // @[Mux.scala 31:69:@39549.4]
  assign _T_94576 = _T_94445 ? 16'h8 : _T_94575; // @[Mux.scala 31:69:@39550.4]
  assign _T_94577 = _T_94442 ? 16'h4 : _T_94576; // @[Mux.scala 31:69:@39551.4]
  assign _T_94578 = _T_94439 ? 16'h2 : _T_94577; // @[Mux.scala 31:69:@39552.4]
  assign _T_94579 = _T_94436 ? 16'h1 : _T_94578; // @[Mux.scala 31:69:@39553.4]
  assign _T_94580 = _T_94579[0]; // @[OneHot.scala 66:30:@39554.4]
  assign _T_94581 = _T_94579[1]; // @[OneHot.scala 66:30:@39555.4]
  assign _T_94582 = _T_94579[2]; // @[OneHot.scala 66:30:@39556.4]
  assign _T_94583 = _T_94579[3]; // @[OneHot.scala 66:30:@39557.4]
  assign _T_94584 = _T_94579[4]; // @[OneHot.scala 66:30:@39558.4]
  assign _T_94585 = _T_94579[5]; // @[OneHot.scala 66:30:@39559.4]
  assign _T_94586 = _T_94579[6]; // @[OneHot.scala 66:30:@39560.4]
  assign _T_94587 = _T_94579[7]; // @[OneHot.scala 66:30:@39561.4]
  assign _T_94588 = _T_94579[8]; // @[OneHot.scala 66:30:@39562.4]
  assign _T_94589 = _T_94579[9]; // @[OneHot.scala 66:30:@39563.4]
  assign _T_94590 = _T_94579[10]; // @[OneHot.scala 66:30:@39564.4]
  assign _T_94591 = _T_94579[11]; // @[OneHot.scala 66:30:@39565.4]
  assign _T_94592 = _T_94579[12]; // @[OneHot.scala 66:30:@39566.4]
  assign _T_94593 = _T_94579[13]; // @[OneHot.scala 66:30:@39567.4]
  assign _T_94594 = _T_94579[14]; // @[OneHot.scala 66:30:@39568.4]
  assign _T_94595 = _T_94579[15]; // @[OneHot.scala 66:30:@39569.4]
  assign _T_94636 = _T_94436 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39587.4]
  assign _T_94637 = _T_94481 ? 16'h4000 : _T_94636; // @[Mux.scala 31:69:@39588.4]
  assign _T_94638 = _T_94478 ? 16'h2000 : _T_94637; // @[Mux.scala 31:69:@39589.4]
  assign _T_94639 = _T_94475 ? 16'h1000 : _T_94638; // @[Mux.scala 31:69:@39590.4]
  assign _T_94640 = _T_94472 ? 16'h800 : _T_94639; // @[Mux.scala 31:69:@39591.4]
  assign _T_94641 = _T_94469 ? 16'h400 : _T_94640; // @[Mux.scala 31:69:@39592.4]
  assign _T_94642 = _T_94466 ? 16'h200 : _T_94641; // @[Mux.scala 31:69:@39593.4]
  assign _T_94643 = _T_94463 ? 16'h100 : _T_94642; // @[Mux.scala 31:69:@39594.4]
  assign _T_94644 = _T_94460 ? 16'h80 : _T_94643; // @[Mux.scala 31:69:@39595.4]
  assign _T_94645 = _T_94457 ? 16'h40 : _T_94644; // @[Mux.scala 31:69:@39596.4]
  assign _T_94646 = _T_94454 ? 16'h20 : _T_94645; // @[Mux.scala 31:69:@39597.4]
  assign _T_94647 = _T_94451 ? 16'h10 : _T_94646; // @[Mux.scala 31:69:@39598.4]
  assign _T_94648 = _T_94448 ? 16'h8 : _T_94647; // @[Mux.scala 31:69:@39599.4]
  assign _T_94649 = _T_94445 ? 16'h4 : _T_94648; // @[Mux.scala 31:69:@39600.4]
  assign _T_94650 = _T_94442 ? 16'h2 : _T_94649; // @[Mux.scala 31:69:@39601.4]
  assign _T_94651 = _T_94439 ? 16'h1 : _T_94650; // @[Mux.scala 31:69:@39602.4]
  assign _T_94652 = _T_94651[0]; // @[OneHot.scala 66:30:@39603.4]
  assign _T_94653 = _T_94651[1]; // @[OneHot.scala 66:30:@39604.4]
  assign _T_94654 = _T_94651[2]; // @[OneHot.scala 66:30:@39605.4]
  assign _T_94655 = _T_94651[3]; // @[OneHot.scala 66:30:@39606.4]
  assign _T_94656 = _T_94651[4]; // @[OneHot.scala 66:30:@39607.4]
  assign _T_94657 = _T_94651[5]; // @[OneHot.scala 66:30:@39608.4]
  assign _T_94658 = _T_94651[6]; // @[OneHot.scala 66:30:@39609.4]
  assign _T_94659 = _T_94651[7]; // @[OneHot.scala 66:30:@39610.4]
  assign _T_94660 = _T_94651[8]; // @[OneHot.scala 66:30:@39611.4]
  assign _T_94661 = _T_94651[9]; // @[OneHot.scala 66:30:@39612.4]
  assign _T_94662 = _T_94651[10]; // @[OneHot.scala 66:30:@39613.4]
  assign _T_94663 = _T_94651[11]; // @[OneHot.scala 66:30:@39614.4]
  assign _T_94664 = _T_94651[12]; // @[OneHot.scala 66:30:@39615.4]
  assign _T_94665 = _T_94651[13]; // @[OneHot.scala 66:30:@39616.4]
  assign _T_94666 = _T_94651[14]; // @[OneHot.scala 66:30:@39617.4]
  assign _T_94667 = _T_94651[15]; // @[OneHot.scala 66:30:@39618.4]
  assign _T_94708 = _T_94439 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39636.4]
  assign _T_94709 = _T_94436 ? 16'h4000 : _T_94708; // @[Mux.scala 31:69:@39637.4]
  assign _T_94710 = _T_94481 ? 16'h2000 : _T_94709; // @[Mux.scala 31:69:@39638.4]
  assign _T_94711 = _T_94478 ? 16'h1000 : _T_94710; // @[Mux.scala 31:69:@39639.4]
  assign _T_94712 = _T_94475 ? 16'h800 : _T_94711; // @[Mux.scala 31:69:@39640.4]
  assign _T_94713 = _T_94472 ? 16'h400 : _T_94712; // @[Mux.scala 31:69:@39641.4]
  assign _T_94714 = _T_94469 ? 16'h200 : _T_94713; // @[Mux.scala 31:69:@39642.4]
  assign _T_94715 = _T_94466 ? 16'h100 : _T_94714; // @[Mux.scala 31:69:@39643.4]
  assign _T_94716 = _T_94463 ? 16'h80 : _T_94715; // @[Mux.scala 31:69:@39644.4]
  assign _T_94717 = _T_94460 ? 16'h40 : _T_94716; // @[Mux.scala 31:69:@39645.4]
  assign _T_94718 = _T_94457 ? 16'h20 : _T_94717; // @[Mux.scala 31:69:@39646.4]
  assign _T_94719 = _T_94454 ? 16'h10 : _T_94718; // @[Mux.scala 31:69:@39647.4]
  assign _T_94720 = _T_94451 ? 16'h8 : _T_94719; // @[Mux.scala 31:69:@39648.4]
  assign _T_94721 = _T_94448 ? 16'h4 : _T_94720; // @[Mux.scala 31:69:@39649.4]
  assign _T_94722 = _T_94445 ? 16'h2 : _T_94721; // @[Mux.scala 31:69:@39650.4]
  assign _T_94723 = _T_94442 ? 16'h1 : _T_94722; // @[Mux.scala 31:69:@39651.4]
  assign _T_94724 = _T_94723[0]; // @[OneHot.scala 66:30:@39652.4]
  assign _T_94725 = _T_94723[1]; // @[OneHot.scala 66:30:@39653.4]
  assign _T_94726 = _T_94723[2]; // @[OneHot.scala 66:30:@39654.4]
  assign _T_94727 = _T_94723[3]; // @[OneHot.scala 66:30:@39655.4]
  assign _T_94728 = _T_94723[4]; // @[OneHot.scala 66:30:@39656.4]
  assign _T_94729 = _T_94723[5]; // @[OneHot.scala 66:30:@39657.4]
  assign _T_94730 = _T_94723[6]; // @[OneHot.scala 66:30:@39658.4]
  assign _T_94731 = _T_94723[7]; // @[OneHot.scala 66:30:@39659.4]
  assign _T_94732 = _T_94723[8]; // @[OneHot.scala 66:30:@39660.4]
  assign _T_94733 = _T_94723[9]; // @[OneHot.scala 66:30:@39661.4]
  assign _T_94734 = _T_94723[10]; // @[OneHot.scala 66:30:@39662.4]
  assign _T_94735 = _T_94723[11]; // @[OneHot.scala 66:30:@39663.4]
  assign _T_94736 = _T_94723[12]; // @[OneHot.scala 66:30:@39664.4]
  assign _T_94737 = _T_94723[13]; // @[OneHot.scala 66:30:@39665.4]
  assign _T_94738 = _T_94723[14]; // @[OneHot.scala 66:30:@39666.4]
  assign _T_94739 = _T_94723[15]; // @[OneHot.scala 66:30:@39667.4]
  assign _T_94780 = _T_94442 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39685.4]
  assign _T_94781 = _T_94439 ? 16'h4000 : _T_94780; // @[Mux.scala 31:69:@39686.4]
  assign _T_94782 = _T_94436 ? 16'h2000 : _T_94781; // @[Mux.scala 31:69:@39687.4]
  assign _T_94783 = _T_94481 ? 16'h1000 : _T_94782; // @[Mux.scala 31:69:@39688.4]
  assign _T_94784 = _T_94478 ? 16'h800 : _T_94783; // @[Mux.scala 31:69:@39689.4]
  assign _T_94785 = _T_94475 ? 16'h400 : _T_94784; // @[Mux.scala 31:69:@39690.4]
  assign _T_94786 = _T_94472 ? 16'h200 : _T_94785; // @[Mux.scala 31:69:@39691.4]
  assign _T_94787 = _T_94469 ? 16'h100 : _T_94786; // @[Mux.scala 31:69:@39692.4]
  assign _T_94788 = _T_94466 ? 16'h80 : _T_94787; // @[Mux.scala 31:69:@39693.4]
  assign _T_94789 = _T_94463 ? 16'h40 : _T_94788; // @[Mux.scala 31:69:@39694.4]
  assign _T_94790 = _T_94460 ? 16'h20 : _T_94789; // @[Mux.scala 31:69:@39695.4]
  assign _T_94791 = _T_94457 ? 16'h10 : _T_94790; // @[Mux.scala 31:69:@39696.4]
  assign _T_94792 = _T_94454 ? 16'h8 : _T_94791; // @[Mux.scala 31:69:@39697.4]
  assign _T_94793 = _T_94451 ? 16'h4 : _T_94792; // @[Mux.scala 31:69:@39698.4]
  assign _T_94794 = _T_94448 ? 16'h2 : _T_94793; // @[Mux.scala 31:69:@39699.4]
  assign _T_94795 = _T_94445 ? 16'h1 : _T_94794; // @[Mux.scala 31:69:@39700.4]
  assign _T_94796 = _T_94795[0]; // @[OneHot.scala 66:30:@39701.4]
  assign _T_94797 = _T_94795[1]; // @[OneHot.scala 66:30:@39702.4]
  assign _T_94798 = _T_94795[2]; // @[OneHot.scala 66:30:@39703.4]
  assign _T_94799 = _T_94795[3]; // @[OneHot.scala 66:30:@39704.4]
  assign _T_94800 = _T_94795[4]; // @[OneHot.scala 66:30:@39705.4]
  assign _T_94801 = _T_94795[5]; // @[OneHot.scala 66:30:@39706.4]
  assign _T_94802 = _T_94795[6]; // @[OneHot.scala 66:30:@39707.4]
  assign _T_94803 = _T_94795[7]; // @[OneHot.scala 66:30:@39708.4]
  assign _T_94804 = _T_94795[8]; // @[OneHot.scala 66:30:@39709.4]
  assign _T_94805 = _T_94795[9]; // @[OneHot.scala 66:30:@39710.4]
  assign _T_94806 = _T_94795[10]; // @[OneHot.scala 66:30:@39711.4]
  assign _T_94807 = _T_94795[11]; // @[OneHot.scala 66:30:@39712.4]
  assign _T_94808 = _T_94795[12]; // @[OneHot.scala 66:30:@39713.4]
  assign _T_94809 = _T_94795[13]; // @[OneHot.scala 66:30:@39714.4]
  assign _T_94810 = _T_94795[14]; // @[OneHot.scala 66:30:@39715.4]
  assign _T_94811 = _T_94795[15]; // @[OneHot.scala 66:30:@39716.4]
  assign _T_94852 = _T_94445 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39734.4]
  assign _T_94853 = _T_94442 ? 16'h4000 : _T_94852; // @[Mux.scala 31:69:@39735.4]
  assign _T_94854 = _T_94439 ? 16'h2000 : _T_94853; // @[Mux.scala 31:69:@39736.4]
  assign _T_94855 = _T_94436 ? 16'h1000 : _T_94854; // @[Mux.scala 31:69:@39737.4]
  assign _T_94856 = _T_94481 ? 16'h800 : _T_94855; // @[Mux.scala 31:69:@39738.4]
  assign _T_94857 = _T_94478 ? 16'h400 : _T_94856; // @[Mux.scala 31:69:@39739.4]
  assign _T_94858 = _T_94475 ? 16'h200 : _T_94857; // @[Mux.scala 31:69:@39740.4]
  assign _T_94859 = _T_94472 ? 16'h100 : _T_94858; // @[Mux.scala 31:69:@39741.4]
  assign _T_94860 = _T_94469 ? 16'h80 : _T_94859; // @[Mux.scala 31:69:@39742.4]
  assign _T_94861 = _T_94466 ? 16'h40 : _T_94860; // @[Mux.scala 31:69:@39743.4]
  assign _T_94862 = _T_94463 ? 16'h20 : _T_94861; // @[Mux.scala 31:69:@39744.4]
  assign _T_94863 = _T_94460 ? 16'h10 : _T_94862; // @[Mux.scala 31:69:@39745.4]
  assign _T_94864 = _T_94457 ? 16'h8 : _T_94863; // @[Mux.scala 31:69:@39746.4]
  assign _T_94865 = _T_94454 ? 16'h4 : _T_94864; // @[Mux.scala 31:69:@39747.4]
  assign _T_94866 = _T_94451 ? 16'h2 : _T_94865; // @[Mux.scala 31:69:@39748.4]
  assign _T_94867 = _T_94448 ? 16'h1 : _T_94866; // @[Mux.scala 31:69:@39749.4]
  assign _T_94868 = _T_94867[0]; // @[OneHot.scala 66:30:@39750.4]
  assign _T_94869 = _T_94867[1]; // @[OneHot.scala 66:30:@39751.4]
  assign _T_94870 = _T_94867[2]; // @[OneHot.scala 66:30:@39752.4]
  assign _T_94871 = _T_94867[3]; // @[OneHot.scala 66:30:@39753.4]
  assign _T_94872 = _T_94867[4]; // @[OneHot.scala 66:30:@39754.4]
  assign _T_94873 = _T_94867[5]; // @[OneHot.scala 66:30:@39755.4]
  assign _T_94874 = _T_94867[6]; // @[OneHot.scala 66:30:@39756.4]
  assign _T_94875 = _T_94867[7]; // @[OneHot.scala 66:30:@39757.4]
  assign _T_94876 = _T_94867[8]; // @[OneHot.scala 66:30:@39758.4]
  assign _T_94877 = _T_94867[9]; // @[OneHot.scala 66:30:@39759.4]
  assign _T_94878 = _T_94867[10]; // @[OneHot.scala 66:30:@39760.4]
  assign _T_94879 = _T_94867[11]; // @[OneHot.scala 66:30:@39761.4]
  assign _T_94880 = _T_94867[12]; // @[OneHot.scala 66:30:@39762.4]
  assign _T_94881 = _T_94867[13]; // @[OneHot.scala 66:30:@39763.4]
  assign _T_94882 = _T_94867[14]; // @[OneHot.scala 66:30:@39764.4]
  assign _T_94883 = _T_94867[15]; // @[OneHot.scala 66:30:@39765.4]
  assign _T_94924 = _T_94448 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39783.4]
  assign _T_94925 = _T_94445 ? 16'h4000 : _T_94924; // @[Mux.scala 31:69:@39784.4]
  assign _T_94926 = _T_94442 ? 16'h2000 : _T_94925; // @[Mux.scala 31:69:@39785.4]
  assign _T_94927 = _T_94439 ? 16'h1000 : _T_94926; // @[Mux.scala 31:69:@39786.4]
  assign _T_94928 = _T_94436 ? 16'h800 : _T_94927; // @[Mux.scala 31:69:@39787.4]
  assign _T_94929 = _T_94481 ? 16'h400 : _T_94928; // @[Mux.scala 31:69:@39788.4]
  assign _T_94930 = _T_94478 ? 16'h200 : _T_94929; // @[Mux.scala 31:69:@39789.4]
  assign _T_94931 = _T_94475 ? 16'h100 : _T_94930; // @[Mux.scala 31:69:@39790.4]
  assign _T_94932 = _T_94472 ? 16'h80 : _T_94931; // @[Mux.scala 31:69:@39791.4]
  assign _T_94933 = _T_94469 ? 16'h40 : _T_94932; // @[Mux.scala 31:69:@39792.4]
  assign _T_94934 = _T_94466 ? 16'h20 : _T_94933; // @[Mux.scala 31:69:@39793.4]
  assign _T_94935 = _T_94463 ? 16'h10 : _T_94934; // @[Mux.scala 31:69:@39794.4]
  assign _T_94936 = _T_94460 ? 16'h8 : _T_94935; // @[Mux.scala 31:69:@39795.4]
  assign _T_94937 = _T_94457 ? 16'h4 : _T_94936; // @[Mux.scala 31:69:@39796.4]
  assign _T_94938 = _T_94454 ? 16'h2 : _T_94937; // @[Mux.scala 31:69:@39797.4]
  assign _T_94939 = _T_94451 ? 16'h1 : _T_94938; // @[Mux.scala 31:69:@39798.4]
  assign _T_94940 = _T_94939[0]; // @[OneHot.scala 66:30:@39799.4]
  assign _T_94941 = _T_94939[1]; // @[OneHot.scala 66:30:@39800.4]
  assign _T_94942 = _T_94939[2]; // @[OneHot.scala 66:30:@39801.4]
  assign _T_94943 = _T_94939[3]; // @[OneHot.scala 66:30:@39802.4]
  assign _T_94944 = _T_94939[4]; // @[OneHot.scala 66:30:@39803.4]
  assign _T_94945 = _T_94939[5]; // @[OneHot.scala 66:30:@39804.4]
  assign _T_94946 = _T_94939[6]; // @[OneHot.scala 66:30:@39805.4]
  assign _T_94947 = _T_94939[7]; // @[OneHot.scala 66:30:@39806.4]
  assign _T_94948 = _T_94939[8]; // @[OneHot.scala 66:30:@39807.4]
  assign _T_94949 = _T_94939[9]; // @[OneHot.scala 66:30:@39808.4]
  assign _T_94950 = _T_94939[10]; // @[OneHot.scala 66:30:@39809.4]
  assign _T_94951 = _T_94939[11]; // @[OneHot.scala 66:30:@39810.4]
  assign _T_94952 = _T_94939[12]; // @[OneHot.scala 66:30:@39811.4]
  assign _T_94953 = _T_94939[13]; // @[OneHot.scala 66:30:@39812.4]
  assign _T_94954 = _T_94939[14]; // @[OneHot.scala 66:30:@39813.4]
  assign _T_94955 = _T_94939[15]; // @[OneHot.scala 66:30:@39814.4]
  assign _T_94996 = _T_94451 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39832.4]
  assign _T_94997 = _T_94448 ? 16'h4000 : _T_94996; // @[Mux.scala 31:69:@39833.4]
  assign _T_94998 = _T_94445 ? 16'h2000 : _T_94997; // @[Mux.scala 31:69:@39834.4]
  assign _T_94999 = _T_94442 ? 16'h1000 : _T_94998; // @[Mux.scala 31:69:@39835.4]
  assign _T_95000 = _T_94439 ? 16'h800 : _T_94999; // @[Mux.scala 31:69:@39836.4]
  assign _T_95001 = _T_94436 ? 16'h400 : _T_95000; // @[Mux.scala 31:69:@39837.4]
  assign _T_95002 = _T_94481 ? 16'h200 : _T_95001; // @[Mux.scala 31:69:@39838.4]
  assign _T_95003 = _T_94478 ? 16'h100 : _T_95002; // @[Mux.scala 31:69:@39839.4]
  assign _T_95004 = _T_94475 ? 16'h80 : _T_95003; // @[Mux.scala 31:69:@39840.4]
  assign _T_95005 = _T_94472 ? 16'h40 : _T_95004; // @[Mux.scala 31:69:@39841.4]
  assign _T_95006 = _T_94469 ? 16'h20 : _T_95005; // @[Mux.scala 31:69:@39842.4]
  assign _T_95007 = _T_94466 ? 16'h10 : _T_95006; // @[Mux.scala 31:69:@39843.4]
  assign _T_95008 = _T_94463 ? 16'h8 : _T_95007; // @[Mux.scala 31:69:@39844.4]
  assign _T_95009 = _T_94460 ? 16'h4 : _T_95008; // @[Mux.scala 31:69:@39845.4]
  assign _T_95010 = _T_94457 ? 16'h2 : _T_95009; // @[Mux.scala 31:69:@39846.4]
  assign _T_95011 = _T_94454 ? 16'h1 : _T_95010; // @[Mux.scala 31:69:@39847.4]
  assign _T_95012 = _T_95011[0]; // @[OneHot.scala 66:30:@39848.4]
  assign _T_95013 = _T_95011[1]; // @[OneHot.scala 66:30:@39849.4]
  assign _T_95014 = _T_95011[2]; // @[OneHot.scala 66:30:@39850.4]
  assign _T_95015 = _T_95011[3]; // @[OneHot.scala 66:30:@39851.4]
  assign _T_95016 = _T_95011[4]; // @[OneHot.scala 66:30:@39852.4]
  assign _T_95017 = _T_95011[5]; // @[OneHot.scala 66:30:@39853.4]
  assign _T_95018 = _T_95011[6]; // @[OneHot.scala 66:30:@39854.4]
  assign _T_95019 = _T_95011[7]; // @[OneHot.scala 66:30:@39855.4]
  assign _T_95020 = _T_95011[8]; // @[OneHot.scala 66:30:@39856.4]
  assign _T_95021 = _T_95011[9]; // @[OneHot.scala 66:30:@39857.4]
  assign _T_95022 = _T_95011[10]; // @[OneHot.scala 66:30:@39858.4]
  assign _T_95023 = _T_95011[11]; // @[OneHot.scala 66:30:@39859.4]
  assign _T_95024 = _T_95011[12]; // @[OneHot.scala 66:30:@39860.4]
  assign _T_95025 = _T_95011[13]; // @[OneHot.scala 66:30:@39861.4]
  assign _T_95026 = _T_95011[14]; // @[OneHot.scala 66:30:@39862.4]
  assign _T_95027 = _T_95011[15]; // @[OneHot.scala 66:30:@39863.4]
  assign _T_95068 = _T_94454 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39881.4]
  assign _T_95069 = _T_94451 ? 16'h4000 : _T_95068; // @[Mux.scala 31:69:@39882.4]
  assign _T_95070 = _T_94448 ? 16'h2000 : _T_95069; // @[Mux.scala 31:69:@39883.4]
  assign _T_95071 = _T_94445 ? 16'h1000 : _T_95070; // @[Mux.scala 31:69:@39884.4]
  assign _T_95072 = _T_94442 ? 16'h800 : _T_95071; // @[Mux.scala 31:69:@39885.4]
  assign _T_95073 = _T_94439 ? 16'h400 : _T_95072; // @[Mux.scala 31:69:@39886.4]
  assign _T_95074 = _T_94436 ? 16'h200 : _T_95073; // @[Mux.scala 31:69:@39887.4]
  assign _T_95075 = _T_94481 ? 16'h100 : _T_95074; // @[Mux.scala 31:69:@39888.4]
  assign _T_95076 = _T_94478 ? 16'h80 : _T_95075; // @[Mux.scala 31:69:@39889.4]
  assign _T_95077 = _T_94475 ? 16'h40 : _T_95076; // @[Mux.scala 31:69:@39890.4]
  assign _T_95078 = _T_94472 ? 16'h20 : _T_95077; // @[Mux.scala 31:69:@39891.4]
  assign _T_95079 = _T_94469 ? 16'h10 : _T_95078; // @[Mux.scala 31:69:@39892.4]
  assign _T_95080 = _T_94466 ? 16'h8 : _T_95079; // @[Mux.scala 31:69:@39893.4]
  assign _T_95081 = _T_94463 ? 16'h4 : _T_95080; // @[Mux.scala 31:69:@39894.4]
  assign _T_95082 = _T_94460 ? 16'h2 : _T_95081; // @[Mux.scala 31:69:@39895.4]
  assign _T_95083 = _T_94457 ? 16'h1 : _T_95082; // @[Mux.scala 31:69:@39896.4]
  assign _T_95084 = _T_95083[0]; // @[OneHot.scala 66:30:@39897.4]
  assign _T_95085 = _T_95083[1]; // @[OneHot.scala 66:30:@39898.4]
  assign _T_95086 = _T_95083[2]; // @[OneHot.scala 66:30:@39899.4]
  assign _T_95087 = _T_95083[3]; // @[OneHot.scala 66:30:@39900.4]
  assign _T_95088 = _T_95083[4]; // @[OneHot.scala 66:30:@39901.4]
  assign _T_95089 = _T_95083[5]; // @[OneHot.scala 66:30:@39902.4]
  assign _T_95090 = _T_95083[6]; // @[OneHot.scala 66:30:@39903.4]
  assign _T_95091 = _T_95083[7]; // @[OneHot.scala 66:30:@39904.4]
  assign _T_95092 = _T_95083[8]; // @[OneHot.scala 66:30:@39905.4]
  assign _T_95093 = _T_95083[9]; // @[OneHot.scala 66:30:@39906.4]
  assign _T_95094 = _T_95083[10]; // @[OneHot.scala 66:30:@39907.4]
  assign _T_95095 = _T_95083[11]; // @[OneHot.scala 66:30:@39908.4]
  assign _T_95096 = _T_95083[12]; // @[OneHot.scala 66:30:@39909.4]
  assign _T_95097 = _T_95083[13]; // @[OneHot.scala 66:30:@39910.4]
  assign _T_95098 = _T_95083[14]; // @[OneHot.scala 66:30:@39911.4]
  assign _T_95099 = _T_95083[15]; // @[OneHot.scala 66:30:@39912.4]
  assign _T_95140 = _T_94457 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39930.4]
  assign _T_95141 = _T_94454 ? 16'h4000 : _T_95140; // @[Mux.scala 31:69:@39931.4]
  assign _T_95142 = _T_94451 ? 16'h2000 : _T_95141; // @[Mux.scala 31:69:@39932.4]
  assign _T_95143 = _T_94448 ? 16'h1000 : _T_95142; // @[Mux.scala 31:69:@39933.4]
  assign _T_95144 = _T_94445 ? 16'h800 : _T_95143; // @[Mux.scala 31:69:@39934.4]
  assign _T_95145 = _T_94442 ? 16'h400 : _T_95144; // @[Mux.scala 31:69:@39935.4]
  assign _T_95146 = _T_94439 ? 16'h200 : _T_95145; // @[Mux.scala 31:69:@39936.4]
  assign _T_95147 = _T_94436 ? 16'h100 : _T_95146; // @[Mux.scala 31:69:@39937.4]
  assign _T_95148 = _T_94481 ? 16'h80 : _T_95147; // @[Mux.scala 31:69:@39938.4]
  assign _T_95149 = _T_94478 ? 16'h40 : _T_95148; // @[Mux.scala 31:69:@39939.4]
  assign _T_95150 = _T_94475 ? 16'h20 : _T_95149; // @[Mux.scala 31:69:@39940.4]
  assign _T_95151 = _T_94472 ? 16'h10 : _T_95150; // @[Mux.scala 31:69:@39941.4]
  assign _T_95152 = _T_94469 ? 16'h8 : _T_95151; // @[Mux.scala 31:69:@39942.4]
  assign _T_95153 = _T_94466 ? 16'h4 : _T_95152; // @[Mux.scala 31:69:@39943.4]
  assign _T_95154 = _T_94463 ? 16'h2 : _T_95153; // @[Mux.scala 31:69:@39944.4]
  assign _T_95155 = _T_94460 ? 16'h1 : _T_95154; // @[Mux.scala 31:69:@39945.4]
  assign _T_95156 = _T_95155[0]; // @[OneHot.scala 66:30:@39946.4]
  assign _T_95157 = _T_95155[1]; // @[OneHot.scala 66:30:@39947.4]
  assign _T_95158 = _T_95155[2]; // @[OneHot.scala 66:30:@39948.4]
  assign _T_95159 = _T_95155[3]; // @[OneHot.scala 66:30:@39949.4]
  assign _T_95160 = _T_95155[4]; // @[OneHot.scala 66:30:@39950.4]
  assign _T_95161 = _T_95155[5]; // @[OneHot.scala 66:30:@39951.4]
  assign _T_95162 = _T_95155[6]; // @[OneHot.scala 66:30:@39952.4]
  assign _T_95163 = _T_95155[7]; // @[OneHot.scala 66:30:@39953.4]
  assign _T_95164 = _T_95155[8]; // @[OneHot.scala 66:30:@39954.4]
  assign _T_95165 = _T_95155[9]; // @[OneHot.scala 66:30:@39955.4]
  assign _T_95166 = _T_95155[10]; // @[OneHot.scala 66:30:@39956.4]
  assign _T_95167 = _T_95155[11]; // @[OneHot.scala 66:30:@39957.4]
  assign _T_95168 = _T_95155[12]; // @[OneHot.scala 66:30:@39958.4]
  assign _T_95169 = _T_95155[13]; // @[OneHot.scala 66:30:@39959.4]
  assign _T_95170 = _T_95155[14]; // @[OneHot.scala 66:30:@39960.4]
  assign _T_95171 = _T_95155[15]; // @[OneHot.scala 66:30:@39961.4]
  assign _T_95212 = _T_94460 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39979.4]
  assign _T_95213 = _T_94457 ? 16'h4000 : _T_95212; // @[Mux.scala 31:69:@39980.4]
  assign _T_95214 = _T_94454 ? 16'h2000 : _T_95213; // @[Mux.scala 31:69:@39981.4]
  assign _T_95215 = _T_94451 ? 16'h1000 : _T_95214; // @[Mux.scala 31:69:@39982.4]
  assign _T_95216 = _T_94448 ? 16'h800 : _T_95215; // @[Mux.scala 31:69:@39983.4]
  assign _T_95217 = _T_94445 ? 16'h400 : _T_95216; // @[Mux.scala 31:69:@39984.4]
  assign _T_95218 = _T_94442 ? 16'h200 : _T_95217; // @[Mux.scala 31:69:@39985.4]
  assign _T_95219 = _T_94439 ? 16'h100 : _T_95218; // @[Mux.scala 31:69:@39986.4]
  assign _T_95220 = _T_94436 ? 16'h80 : _T_95219; // @[Mux.scala 31:69:@39987.4]
  assign _T_95221 = _T_94481 ? 16'h40 : _T_95220; // @[Mux.scala 31:69:@39988.4]
  assign _T_95222 = _T_94478 ? 16'h20 : _T_95221; // @[Mux.scala 31:69:@39989.4]
  assign _T_95223 = _T_94475 ? 16'h10 : _T_95222; // @[Mux.scala 31:69:@39990.4]
  assign _T_95224 = _T_94472 ? 16'h8 : _T_95223; // @[Mux.scala 31:69:@39991.4]
  assign _T_95225 = _T_94469 ? 16'h4 : _T_95224; // @[Mux.scala 31:69:@39992.4]
  assign _T_95226 = _T_94466 ? 16'h2 : _T_95225; // @[Mux.scala 31:69:@39993.4]
  assign _T_95227 = _T_94463 ? 16'h1 : _T_95226; // @[Mux.scala 31:69:@39994.4]
  assign _T_95228 = _T_95227[0]; // @[OneHot.scala 66:30:@39995.4]
  assign _T_95229 = _T_95227[1]; // @[OneHot.scala 66:30:@39996.4]
  assign _T_95230 = _T_95227[2]; // @[OneHot.scala 66:30:@39997.4]
  assign _T_95231 = _T_95227[3]; // @[OneHot.scala 66:30:@39998.4]
  assign _T_95232 = _T_95227[4]; // @[OneHot.scala 66:30:@39999.4]
  assign _T_95233 = _T_95227[5]; // @[OneHot.scala 66:30:@40000.4]
  assign _T_95234 = _T_95227[6]; // @[OneHot.scala 66:30:@40001.4]
  assign _T_95235 = _T_95227[7]; // @[OneHot.scala 66:30:@40002.4]
  assign _T_95236 = _T_95227[8]; // @[OneHot.scala 66:30:@40003.4]
  assign _T_95237 = _T_95227[9]; // @[OneHot.scala 66:30:@40004.4]
  assign _T_95238 = _T_95227[10]; // @[OneHot.scala 66:30:@40005.4]
  assign _T_95239 = _T_95227[11]; // @[OneHot.scala 66:30:@40006.4]
  assign _T_95240 = _T_95227[12]; // @[OneHot.scala 66:30:@40007.4]
  assign _T_95241 = _T_95227[13]; // @[OneHot.scala 66:30:@40008.4]
  assign _T_95242 = _T_95227[14]; // @[OneHot.scala 66:30:@40009.4]
  assign _T_95243 = _T_95227[15]; // @[OneHot.scala 66:30:@40010.4]
  assign _T_95284 = _T_94463 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40028.4]
  assign _T_95285 = _T_94460 ? 16'h4000 : _T_95284; // @[Mux.scala 31:69:@40029.4]
  assign _T_95286 = _T_94457 ? 16'h2000 : _T_95285; // @[Mux.scala 31:69:@40030.4]
  assign _T_95287 = _T_94454 ? 16'h1000 : _T_95286; // @[Mux.scala 31:69:@40031.4]
  assign _T_95288 = _T_94451 ? 16'h800 : _T_95287; // @[Mux.scala 31:69:@40032.4]
  assign _T_95289 = _T_94448 ? 16'h400 : _T_95288; // @[Mux.scala 31:69:@40033.4]
  assign _T_95290 = _T_94445 ? 16'h200 : _T_95289; // @[Mux.scala 31:69:@40034.4]
  assign _T_95291 = _T_94442 ? 16'h100 : _T_95290; // @[Mux.scala 31:69:@40035.4]
  assign _T_95292 = _T_94439 ? 16'h80 : _T_95291; // @[Mux.scala 31:69:@40036.4]
  assign _T_95293 = _T_94436 ? 16'h40 : _T_95292; // @[Mux.scala 31:69:@40037.4]
  assign _T_95294 = _T_94481 ? 16'h20 : _T_95293; // @[Mux.scala 31:69:@40038.4]
  assign _T_95295 = _T_94478 ? 16'h10 : _T_95294; // @[Mux.scala 31:69:@40039.4]
  assign _T_95296 = _T_94475 ? 16'h8 : _T_95295; // @[Mux.scala 31:69:@40040.4]
  assign _T_95297 = _T_94472 ? 16'h4 : _T_95296; // @[Mux.scala 31:69:@40041.4]
  assign _T_95298 = _T_94469 ? 16'h2 : _T_95297; // @[Mux.scala 31:69:@40042.4]
  assign _T_95299 = _T_94466 ? 16'h1 : _T_95298; // @[Mux.scala 31:69:@40043.4]
  assign _T_95300 = _T_95299[0]; // @[OneHot.scala 66:30:@40044.4]
  assign _T_95301 = _T_95299[1]; // @[OneHot.scala 66:30:@40045.4]
  assign _T_95302 = _T_95299[2]; // @[OneHot.scala 66:30:@40046.4]
  assign _T_95303 = _T_95299[3]; // @[OneHot.scala 66:30:@40047.4]
  assign _T_95304 = _T_95299[4]; // @[OneHot.scala 66:30:@40048.4]
  assign _T_95305 = _T_95299[5]; // @[OneHot.scala 66:30:@40049.4]
  assign _T_95306 = _T_95299[6]; // @[OneHot.scala 66:30:@40050.4]
  assign _T_95307 = _T_95299[7]; // @[OneHot.scala 66:30:@40051.4]
  assign _T_95308 = _T_95299[8]; // @[OneHot.scala 66:30:@40052.4]
  assign _T_95309 = _T_95299[9]; // @[OneHot.scala 66:30:@40053.4]
  assign _T_95310 = _T_95299[10]; // @[OneHot.scala 66:30:@40054.4]
  assign _T_95311 = _T_95299[11]; // @[OneHot.scala 66:30:@40055.4]
  assign _T_95312 = _T_95299[12]; // @[OneHot.scala 66:30:@40056.4]
  assign _T_95313 = _T_95299[13]; // @[OneHot.scala 66:30:@40057.4]
  assign _T_95314 = _T_95299[14]; // @[OneHot.scala 66:30:@40058.4]
  assign _T_95315 = _T_95299[15]; // @[OneHot.scala 66:30:@40059.4]
  assign _T_95356 = _T_94466 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40077.4]
  assign _T_95357 = _T_94463 ? 16'h4000 : _T_95356; // @[Mux.scala 31:69:@40078.4]
  assign _T_95358 = _T_94460 ? 16'h2000 : _T_95357; // @[Mux.scala 31:69:@40079.4]
  assign _T_95359 = _T_94457 ? 16'h1000 : _T_95358; // @[Mux.scala 31:69:@40080.4]
  assign _T_95360 = _T_94454 ? 16'h800 : _T_95359; // @[Mux.scala 31:69:@40081.4]
  assign _T_95361 = _T_94451 ? 16'h400 : _T_95360; // @[Mux.scala 31:69:@40082.4]
  assign _T_95362 = _T_94448 ? 16'h200 : _T_95361; // @[Mux.scala 31:69:@40083.4]
  assign _T_95363 = _T_94445 ? 16'h100 : _T_95362; // @[Mux.scala 31:69:@40084.4]
  assign _T_95364 = _T_94442 ? 16'h80 : _T_95363; // @[Mux.scala 31:69:@40085.4]
  assign _T_95365 = _T_94439 ? 16'h40 : _T_95364; // @[Mux.scala 31:69:@40086.4]
  assign _T_95366 = _T_94436 ? 16'h20 : _T_95365; // @[Mux.scala 31:69:@40087.4]
  assign _T_95367 = _T_94481 ? 16'h10 : _T_95366; // @[Mux.scala 31:69:@40088.4]
  assign _T_95368 = _T_94478 ? 16'h8 : _T_95367; // @[Mux.scala 31:69:@40089.4]
  assign _T_95369 = _T_94475 ? 16'h4 : _T_95368; // @[Mux.scala 31:69:@40090.4]
  assign _T_95370 = _T_94472 ? 16'h2 : _T_95369; // @[Mux.scala 31:69:@40091.4]
  assign _T_95371 = _T_94469 ? 16'h1 : _T_95370; // @[Mux.scala 31:69:@40092.4]
  assign _T_95372 = _T_95371[0]; // @[OneHot.scala 66:30:@40093.4]
  assign _T_95373 = _T_95371[1]; // @[OneHot.scala 66:30:@40094.4]
  assign _T_95374 = _T_95371[2]; // @[OneHot.scala 66:30:@40095.4]
  assign _T_95375 = _T_95371[3]; // @[OneHot.scala 66:30:@40096.4]
  assign _T_95376 = _T_95371[4]; // @[OneHot.scala 66:30:@40097.4]
  assign _T_95377 = _T_95371[5]; // @[OneHot.scala 66:30:@40098.4]
  assign _T_95378 = _T_95371[6]; // @[OneHot.scala 66:30:@40099.4]
  assign _T_95379 = _T_95371[7]; // @[OneHot.scala 66:30:@40100.4]
  assign _T_95380 = _T_95371[8]; // @[OneHot.scala 66:30:@40101.4]
  assign _T_95381 = _T_95371[9]; // @[OneHot.scala 66:30:@40102.4]
  assign _T_95382 = _T_95371[10]; // @[OneHot.scala 66:30:@40103.4]
  assign _T_95383 = _T_95371[11]; // @[OneHot.scala 66:30:@40104.4]
  assign _T_95384 = _T_95371[12]; // @[OneHot.scala 66:30:@40105.4]
  assign _T_95385 = _T_95371[13]; // @[OneHot.scala 66:30:@40106.4]
  assign _T_95386 = _T_95371[14]; // @[OneHot.scala 66:30:@40107.4]
  assign _T_95387 = _T_95371[15]; // @[OneHot.scala 66:30:@40108.4]
  assign _T_95428 = _T_94469 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40126.4]
  assign _T_95429 = _T_94466 ? 16'h4000 : _T_95428; // @[Mux.scala 31:69:@40127.4]
  assign _T_95430 = _T_94463 ? 16'h2000 : _T_95429; // @[Mux.scala 31:69:@40128.4]
  assign _T_95431 = _T_94460 ? 16'h1000 : _T_95430; // @[Mux.scala 31:69:@40129.4]
  assign _T_95432 = _T_94457 ? 16'h800 : _T_95431; // @[Mux.scala 31:69:@40130.4]
  assign _T_95433 = _T_94454 ? 16'h400 : _T_95432; // @[Mux.scala 31:69:@40131.4]
  assign _T_95434 = _T_94451 ? 16'h200 : _T_95433; // @[Mux.scala 31:69:@40132.4]
  assign _T_95435 = _T_94448 ? 16'h100 : _T_95434; // @[Mux.scala 31:69:@40133.4]
  assign _T_95436 = _T_94445 ? 16'h80 : _T_95435; // @[Mux.scala 31:69:@40134.4]
  assign _T_95437 = _T_94442 ? 16'h40 : _T_95436; // @[Mux.scala 31:69:@40135.4]
  assign _T_95438 = _T_94439 ? 16'h20 : _T_95437; // @[Mux.scala 31:69:@40136.4]
  assign _T_95439 = _T_94436 ? 16'h10 : _T_95438; // @[Mux.scala 31:69:@40137.4]
  assign _T_95440 = _T_94481 ? 16'h8 : _T_95439; // @[Mux.scala 31:69:@40138.4]
  assign _T_95441 = _T_94478 ? 16'h4 : _T_95440; // @[Mux.scala 31:69:@40139.4]
  assign _T_95442 = _T_94475 ? 16'h2 : _T_95441; // @[Mux.scala 31:69:@40140.4]
  assign _T_95443 = _T_94472 ? 16'h1 : _T_95442; // @[Mux.scala 31:69:@40141.4]
  assign _T_95444 = _T_95443[0]; // @[OneHot.scala 66:30:@40142.4]
  assign _T_95445 = _T_95443[1]; // @[OneHot.scala 66:30:@40143.4]
  assign _T_95446 = _T_95443[2]; // @[OneHot.scala 66:30:@40144.4]
  assign _T_95447 = _T_95443[3]; // @[OneHot.scala 66:30:@40145.4]
  assign _T_95448 = _T_95443[4]; // @[OneHot.scala 66:30:@40146.4]
  assign _T_95449 = _T_95443[5]; // @[OneHot.scala 66:30:@40147.4]
  assign _T_95450 = _T_95443[6]; // @[OneHot.scala 66:30:@40148.4]
  assign _T_95451 = _T_95443[7]; // @[OneHot.scala 66:30:@40149.4]
  assign _T_95452 = _T_95443[8]; // @[OneHot.scala 66:30:@40150.4]
  assign _T_95453 = _T_95443[9]; // @[OneHot.scala 66:30:@40151.4]
  assign _T_95454 = _T_95443[10]; // @[OneHot.scala 66:30:@40152.4]
  assign _T_95455 = _T_95443[11]; // @[OneHot.scala 66:30:@40153.4]
  assign _T_95456 = _T_95443[12]; // @[OneHot.scala 66:30:@40154.4]
  assign _T_95457 = _T_95443[13]; // @[OneHot.scala 66:30:@40155.4]
  assign _T_95458 = _T_95443[14]; // @[OneHot.scala 66:30:@40156.4]
  assign _T_95459 = _T_95443[15]; // @[OneHot.scala 66:30:@40157.4]
  assign _T_95500 = _T_94472 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40175.4]
  assign _T_95501 = _T_94469 ? 16'h4000 : _T_95500; // @[Mux.scala 31:69:@40176.4]
  assign _T_95502 = _T_94466 ? 16'h2000 : _T_95501; // @[Mux.scala 31:69:@40177.4]
  assign _T_95503 = _T_94463 ? 16'h1000 : _T_95502; // @[Mux.scala 31:69:@40178.4]
  assign _T_95504 = _T_94460 ? 16'h800 : _T_95503; // @[Mux.scala 31:69:@40179.4]
  assign _T_95505 = _T_94457 ? 16'h400 : _T_95504; // @[Mux.scala 31:69:@40180.4]
  assign _T_95506 = _T_94454 ? 16'h200 : _T_95505; // @[Mux.scala 31:69:@40181.4]
  assign _T_95507 = _T_94451 ? 16'h100 : _T_95506; // @[Mux.scala 31:69:@40182.4]
  assign _T_95508 = _T_94448 ? 16'h80 : _T_95507; // @[Mux.scala 31:69:@40183.4]
  assign _T_95509 = _T_94445 ? 16'h40 : _T_95508; // @[Mux.scala 31:69:@40184.4]
  assign _T_95510 = _T_94442 ? 16'h20 : _T_95509; // @[Mux.scala 31:69:@40185.4]
  assign _T_95511 = _T_94439 ? 16'h10 : _T_95510; // @[Mux.scala 31:69:@40186.4]
  assign _T_95512 = _T_94436 ? 16'h8 : _T_95511; // @[Mux.scala 31:69:@40187.4]
  assign _T_95513 = _T_94481 ? 16'h4 : _T_95512; // @[Mux.scala 31:69:@40188.4]
  assign _T_95514 = _T_94478 ? 16'h2 : _T_95513; // @[Mux.scala 31:69:@40189.4]
  assign _T_95515 = _T_94475 ? 16'h1 : _T_95514; // @[Mux.scala 31:69:@40190.4]
  assign _T_95516 = _T_95515[0]; // @[OneHot.scala 66:30:@40191.4]
  assign _T_95517 = _T_95515[1]; // @[OneHot.scala 66:30:@40192.4]
  assign _T_95518 = _T_95515[2]; // @[OneHot.scala 66:30:@40193.4]
  assign _T_95519 = _T_95515[3]; // @[OneHot.scala 66:30:@40194.4]
  assign _T_95520 = _T_95515[4]; // @[OneHot.scala 66:30:@40195.4]
  assign _T_95521 = _T_95515[5]; // @[OneHot.scala 66:30:@40196.4]
  assign _T_95522 = _T_95515[6]; // @[OneHot.scala 66:30:@40197.4]
  assign _T_95523 = _T_95515[7]; // @[OneHot.scala 66:30:@40198.4]
  assign _T_95524 = _T_95515[8]; // @[OneHot.scala 66:30:@40199.4]
  assign _T_95525 = _T_95515[9]; // @[OneHot.scala 66:30:@40200.4]
  assign _T_95526 = _T_95515[10]; // @[OneHot.scala 66:30:@40201.4]
  assign _T_95527 = _T_95515[11]; // @[OneHot.scala 66:30:@40202.4]
  assign _T_95528 = _T_95515[12]; // @[OneHot.scala 66:30:@40203.4]
  assign _T_95529 = _T_95515[13]; // @[OneHot.scala 66:30:@40204.4]
  assign _T_95530 = _T_95515[14]; // @[OneHot.scala 66:30:@40205.4]
  assign _T_95531 = _T_95515[15]; // @[OneHot.scala 66:30:@40206.4]
  assign _T_95572 = _T_94475 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40224.4]
  assign _T_95573 = _T_94472 ? 16'h4000 : _T_95572; // @[Mux.scala 31:69:@40225.4]
  assign _T_95574 = _T_94469 ? 16'h2000 : _T_95573; // @[Mux.scala 31:69:@40226.4]
  assign _T_95575 = _T_94466 ? 16'h1000 : _T_95574; // @[Mux.scala 31:69:@40227.4]
  assign _T_95576 = _T_94463 ? 16'h800 : _T_95575; // @[Mux.scala 31:69:@40228.4]
  assign _T_95577 = _T_94460 ? 16'h400 : _T_95576; // @[Mux.scala 31:69:@40229.4]
  assign _T_95578 = _T_94457 ? 16'h200 : _T_95577; // @[Mux.scala 31:69:@40230.4]
  assign _T_95579 = _T_94454 ? 16'h100 : _T_95578; // @[Mux.scala 31:69:@40231.4]
  assign _T_95580 = _T_94451 ? 16'h80 : _T_95579; // @[Mux.scala 31:69:@40232.4]
  assign _T_95581 = _T_94448 ? 16'h40 : _T_95580; // @[Mux.scala 31:69:@40233.4]
  assign _T_95582 = _T_94445 ? 16'h20 : _T_95581; // @[Mux.scala 31:69:@40234.4]
  assign _T_95583 = _T_94442 ? 16'h10 : _T_95582; // @[Mux.scala 31:69:@40235.4]
  assign _T_95584 = _T_94439 ? 16'h8 : _T_95583; // @[Mux.scala 31:69:@40236.4]
  assign _T_95585 = _T_94436 ? 16'h4 : _T_95584; // @[Mux.scala 31:69:@40237.4]
  assign _T_95586 = _T_94481 ? 16'h2 : _T_95585; // @[Mux.scala 31:69:@40238.4]
  assign _T_95587 = _T_94478 ? 16'h1 : _T_95586; // @[Mux.scala 31:69:@40239.4]
  assign _T_95588 = _T_95587[0]; // @[OneHot.scala 66:30:@40240.4]
  assign _T_95589 = _T_95587[1]; // @[OneHot.scala 66:30:@40241.4]
  assign _T_95590 = _T_95587[2]; // @[OneHot.scala 66:30:@40242.4]
  assign _T_95591 = _T_95587[3]; // @[OneHot.scala 66:30:@40243.4]
  assign _T_95592 = _T_95587[4]; // @[OneHot.scala 66:30:@40244.4]
  assign _T_95593 = _T_95587[5]; // @[OneHot.scala 66:30:@40245.4]
  assign _T_95594 = _T_95587[6]; // @[OneHot.scala 66:30:@40246.4]
  assign _T_95595 = _T_95587[7]; // @[OneHot.scala 66:30:@40247.4]
  assign _T_95596 = _T_95587[8]; // @[OneHot.scala 66:30:@40248.4]
  assign _T_95597 = _T_95587[9]; // @[OneHot.scala 66:30:@40249.4]
  assign _T_95598 = _T_95587[10]; // @[OneHot.scala 66:30:@40250.4]
  assign _T_95599 = _T_95587[11]; // @[OneHot.scala 66:30:@40251.4]
  assign _T_95600 = _T_95587[12]; // @[OneHot.scala 66:30:@40252.4]
  assign _T_95601 = _T_95587[13]; // @[OneHot.scala 66:30:@40253.4]
  assign _T_95602 = _T_95587[14]; // @[OneHot.scala 66:30:@40254.4]
  assign _T_95603 = _T_95587[15]; // @[OneHot.scala 66:30:@40255.4]
  assign _T_95644 = _T_94478 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40273.4]
  assign _T_95645 = _T_94475 ? 16'h4000 : _T_95644; // @[Mux.scala 31:69:@40274.4]
  assign _T_95646 = _T_94472 ? 16'h2000 : _T_95645; // @[Mux.scala 31:69:@40275.4]
  assign _T_95647 = _T_94469 ? 16'h1000 : _T_95646; // @[Mux.scala 31:69:@40276.4]
  assign _T_95648 = _T_94466 ? 16'h800 : _T_95647; // @[Mux.scala 31:69:@40277.4]
  assign _T_95649 = _T_94463 ? 16'h400 : _T_95648; // @[Mux.scala 31:69:@40278.4]
  assign _T_95650 = _T_94460 ? 16'h200 : _T_95649; // @[Mux.scala 31:69:@40279.4]
  assign _T_95651 = _T_94457 ? 16'h100 : _T_95650; // @[Mux.scala 31:69:@40280.4]
  assign _T_95652 = _T_94454 ? 16'h80 : _T_95651; // @[Mux.scala 31:69:@40281.4]
  assign _T_95653 = _T_94451 ? 16'h40 : _T_95652; // @[Mux.scala 31:69:@40282.4]
  assign _T_95654 = _T_94448 ? 16'h20 : _T_95653; // @[Mux.scala 31:69:@40283.4]
  assign _T_95655 = _T_94445 ? 16'h10 : _T_95654; // @[Mux.scala 31:69:@40284.4]
  assign _T_95656 = _T_94442 ? 16'h8 : _T_95655; // @[Mux.scala 31:69:@40285.4]
  assign _T_95657 = _T_94439 ? 16'h4 : _T_95656; // @[Mux.scala 31:69:@40286.4]
  assign _T_95658 = _T_94436 ? 16'h2 : _T_95657; // @[Mux.scala 31:69:@40287.4]
  assign _T_95659 = _T_94481 ? 16'h1 : _T_95658; // @[Mux.scala 31:69:@40288.4]
  assign _T_95660 = _T_95659[0]; // @[OneHot.scala 66:30:@40289.4]
  assign _T_95661 = _T_95659[1]; // @[OneHot.scala 66:30:@40290.4]
  assign _T_95662 = _T_95659[2]; // @[OneHot.scala 66:30:@40291.4]
  assign _T_95663 = _T_95659[3]; // @[OneHot.scala 66:30:@40292.4]
  assign _T_95664 = _T_95659[4]; // @[OneHot.scala 66:30:@40293.4]
  assign _T_95665 = _T_95659[5]; // @[OneHot.scala 66:30:@40294.4]
  assign _T_95666 = _T_95659[6]; // @[OneHot.scala 66:30:@40295.4]
  assign _T_95667 = _T_95659[7]; // @[OneHot.scala 66:30:@40296.4]
  assign _T_95668 = _T_95659[8]; // @[OneHot.scala 66:30:@40297.4]
  assign _T_95669 = _T_95659[9]; // @[OneHot.scala 66:30:@40298.4]
  assign _T_95670 = _T_95659[10]; // @[OneHot.scala 66:30:@40299.4]
  assign _T_95671 = _T_95659[11]; // @[OneHot.scala 66:30:@40300.4]
  assign _T_95672 = _T_95659[12]; // @[OneHot.scala 66:30:@40301.4]
  assign _T_95673 = _T_95659[13]; // @[OneHot.scala 66:30:@40302.4]
  assign _T_95674 = _T_95659[14]; // @[OneHot.scala 66:30:@40303.4]
  assign _T_95675 = _T_95659[15]; // @[OneHot.scala 66:30:@40304.4]
  assign _T_95740 = {_T_94587,_T_94586,_T_94585,_T_94584,_T_94583,_T_94582,_T_94581,_T_94580}; // @[Mux.scala 19:72:@40328.4]
  assign _T_95748 = {_T_94595,_T_94594,_T_94593,_T_94592,_T_94591,_T_94590,_T_94589,_T_94588,_T_95740}; // @[Mux.scala 19:72:@40336.4]
  assign _T_95750 = _T_90408 ? _T_95748 : 16'h0; // @[Mux.scala 19:72:@40337.4]
  assign _T_95757 = {_T_94658,_T_94657,_T_94656,_T_94655,_T_94654,_T_94653,_T_94652,_T_94667}; // @[Mux.scala 19:72:@40344.4]
  assign _T_95765 = {_T_94666,_T_94665,_T_94664,_T_94663,_T_94662,_T_94661,_T_94660,_T_94659,_T_95757}; // @[Mux.scala 19:72:@40352.4]
  assign _T_95767 = _T_90409 ? _T_95765 : 16'h0; // @[Mux.scala 19:72:@40353.4]
  assign _T_95774 = {_T_94729,_T_94728,_T_94727,_T_94726,_T_94725,_T_94724,_T_94739,_T_94738}; // @[Mux.scala 19:72:@40360.4]
  assign _T_95782 = {_T_94737,_T_94736,_T_94735,_T_94734,_T_94733,_T_94732,_T_94731,_T_94730,_T_95774}; // @[Mux.scala 19:72:@40368.4]
  assign _T_95784 = _T_90410 ? _T_95782 : 16'h0; // @[Mux.scala 19:72:@40369.4]
  assign _T_95791 = {_T_94800,_T_94799,_T_94798,_T_94797,_T_94796,_T_94811,_T_94810,_T_94809}; // @[Mux.scala 19:72:@40376.4]
  assign _T_95799 = {_T_94808,_T_94807,_T_94806,_T_94805,_T_94804,_T_94803,_T_94802,_T_94801,_T_95791}; // @[Mux.scala 19:72:@40384.4]
  assign _T_95801 = _T_90411 ? _T_95799 : 16'h0; // @[Mux.scala 19:72:@40385.4]
  assign _T_95808 = {_T_94871,_T_94870,_T_94869,_T_94868,_T_94883,_T_94882,_T_94881,_T_94880}; // @[Mux.scala 19:72:@40392.4]
  assign _T_95816 = {_T_94879,_T_94878,_T_94877,_T_94876,_T_94875,_T_94874,_T_94873,_T_94872,_T_95808}; // @[Mux.scala 19:72:@40400.4]
  assign _T_95818 = _T_90412 ? _T_95816 : 16'h0; // @[Mux.scala 19:72:@40401.4]
  assign _T_95825 = {_T_94942,_T_94941,_T_94940,_T_94955,_T_94954,_T_94953,_T_94952,_T_94951}; // @[Mux.scala 19:72:@40408.4]
  assign _T_95833 = {_T_94950,_T_94949,_T_94948,_T_94947,_T_94946,_T_94945,_T_94944,_T_94943,_T_95825}; // @[Mux.scala 19:72:@40416.4]
  assign _T_95835 = _T_90413 ? _T_95833 : 16'h0; // @[Mux.scala 19:72:@40417.4]
  assign _T_95842 = {_T_95013,_T_95012,_T_95027,_T_95026,_T_95025,_T_95024,_T_95023,_T_95022}; // @[Mux.scala 19:72:@40424.4]
  assign _T_95850 = {_T_95021,_T_95020,_T_95019,_T_95018,_T_95017,_T_95016,_T_95015,_T_95014,_T_95842}; // @[Mux.scala 19:72:@40432.4]
  assign _T_95852 = _T_90414 ? _T_95850 : 16'h0; // @[Mux.scala 19:72:@40433.4]
  assign _T_95859 = {_T_95084,_T_95099,_T_95098,_T_95097,_T_95096,_T_95095,_T_95094,_T_95093}; // @[Mux.scala 19:72:@40440.4]
  assign _T_95867 = {_T_95092,_T_95091,_T_95090,_T_95089,_T_95088,_T_95087,_T_95086,_T_95085,_T_95859}; // @[Mux.scala 19:72:@40448.4]
  assign _T_95869 = _T_90415 ? _T_95867 : 16'h0; // @[Mux.scala 19:72:@40449.4]
  assign _T_95876 = {_T_95171,_T_95170,_T_95169,_T_95168,_T_95167,_T_95166,_T_95165,_T_95164}; // @[Mux.scala 19:72:@40456.4]
  assign _T_95884 = {_T_95163,_T_95162,_T_95161,_T_95160,_T_95159,_T_95158,_T_95157,_T_95156,_T_95876}; // @[Mux.scala 19:72:@40464.4]
  assign _T_95886 = _T_90416 ? _T_95884 : 16'h0; // @[Mux.scala 19:72:@40465.4]
  assign _T_95893 = {_T_95242,_T_95241,_T_95240,_T_95239,_T_95238,_T_95237,_T_95236,_T_95235}; // @[Mux.scala 19:72:@40472.4]
  assign _T_95901 = {_T_95234,_T_95233,_T_95232,_T_95231,_T_95230,_T_95229,_T_95228,_T_95243,_T_95893}; // @[Mux.scala 19:72:@40480.4]
  assign _T_95903 = _T_90417 ? _T_95901 : 16'h0; // @[Mux.scala 19:72:@40481.4]
  assign _T_95910 = {_T_95313,_T_95312,_T_95311,_T_95310,_T_95309,_T_95308,_T_95307,_T_95306}; // @[Mux.scala 19:72:@40488.4]
  assign _T_95918 = {_T_95305,_T_95304,_T_95303,_T_95302,_T_95301,_T_95300,_T_95315,_T_95314,_T_95910}; // @[Mux.scala 19:72:@40496.4]
  assign _T_95920 = _T_90418 ? _T_95918 : 16'h0; // @[Mux.scala 19:72:@40497.4]
  assign _T_95927 = {_T_95384,_T_95383,_T_95382,_T_95381,_T_95380,_T_95379,_T_95378,_T_95377}; // @[Mux.scala 19:72:@40504.4]
  assign _T_95935 = {_T_95376,_T_95375,_T_95374,_T_95373,_T_95372,_T_95387,_T_95386,_T_95385,_T_95927}; // @[Mux.scala 19:72:@40512.4]
  assign _T_95937 = _T_90419 ? _T_95935 : 16'h0; // @[Mux.scala 19:72:@40513.4]
  assign _T_95944 = {_T_95455,_T_95454,_T_95453,_T_95452,_T_95451,_T_95450,_T_95449,_T_95448}; // @[Mux.scala 19:72:@40520.4]
  assign _T_95952 = {_T_95447,_T_95446,_T_95445,_T_95444,_T_95459,_T_95458,_T_95457,_T_95456,_T_95944}; // @[Mux.scala 19:72:@40528.4]
  assign _T_95954 = _T_90420 ? _T_95952 : 16'h0; // @[Mux.scala 19:72:@40529.4]
  assign _T_95961 = {_T_95526,_T_95525,_T_95524,_T_95523,_T_95522,_T_95521,_T_95520,_T_95519}; // @[Mux.scala 19:72:@40536.4]
  assign _T_95969 = {_T_95518,_T_95517,_T_95516,_T_95531,_T_95530,_T_95529,_T_95528,_T_95527,_T_95961}; // @[Mux.scala 19:72:@40544.4]
  assign _T_95971 = _T_90421 ? _T_95969 : 16'h0; // @[Mux.scala 19:72:@40545.4]
  assign _T_95978 = {_T_95597,_T_95596,_T_95595,_T_95594,_T_95593,_T_95592,_T_95591,_T_95590}; // @[Mux.scala 19:72:@40552.4]
  assign _T_95986 = {_T_95589,_T_95588,_T_95603,_T_95602,_T_95601,_T_95600,_T_95599,_T_95598,_T_95978}; // @[Mux.scala 19:72:@40560.4]
  assign _T_95988 = _T_90422 ? _T_95986 : 16'h0; // @[Mux.scala 19:72:@40561.4]
  assign _T_95995 = {_T_95668,_T_95667,_T_95666,_T_95665,_T_95664,_T_95663,_T_95662,_T_95661}; // @[Mux.scala 19:72:@40568.4]
  assign _T_96003 = {_T_95660,_T_95675,_T_95674,_T_95673,_T_95672,_T_95671,_T_95670,_T_95669,_T_95995}; // @[Mux.scala 19:72:@40576.4]
  assign _T_96005 = _T_90423 ? _T_96003 : 16'h0; // @[Mux.scala 19:72:@40577.4]
  assign _T_96006 = _T_95750 | _T_95767; // @[Mux.scala 19:72:@40578.4]
  assign _T_96007 = _T_96006 | _T_95784; // @[Mux.scala 19:72:@40579.4]
  assign _T_96008 = _T_96007 | _T_95801; // @[Mux.scala 19:72:@40580.4]
  assign _T_96009 = _T_96008 | _T_95818; // @[Mux.scala 19:72:@40581.4]
  assign _T_96010 = _T_96009 | _T_95835; // @[Mux.scala 19:72:@40582.4]
  assign _T_96011 = _T_96010 | _T_95852; // @[Mux.scala 19:72:@40583.4]
  assign _T_96012 = _T_96011 | _T_95869; // @[Mux.scala 19:72:@40584.4]
  assign _T_96013 = _T_96012 | _T_95886; // @[Mux.scala 19:72:@40585.4]
  assign _T_96014 = _T_96013 | _T_95903; // @[Mux.scala 19:72:@40586.4]
  assign _T_96015 = _T_96014 | _T_95920; // @[Mux.scala 19:72:@40587.4]
  assign _T_96016 = _T_96015 | _T_95937; // @[Mux.scala 19:72:@40588.4]
  assign _T_96017 = _T_96016 | _T_95954; // @[Mux.scala 19:72:@40589.4]
  assign _T_96018 = _T_96017 | _T_95971; // @[Mux.scala 19:72:@40590.4]
  assign _T_96019 = _T_96018 | _T_95988; // @[Mux.scala 19:72:@40591.4]
  assign _T_96020 = _T_96019 | _T_96005; // @[Mux.scala 19:72:@40592.4]
  assign inputPriorityPorts_0_0 = _T_96020[0]; // @[Mux.scala 19:72:@40596.4]
  assign inputPriorityPorts_0_1 = _T_96020[1]; // @[Mux.scala 19:72:@40598.4]
  assign inputPriorityPorts_0_2 = _T_96020[2]; // @[Mux.scala 19:72:@40600.4]
  assign inputPriorityPorts_0_3 = _T_96020[3]; // @[Mux.scala 19:72:@40602.4]
  assign inputPriorityPorts_0_4 = _T_96020[4]; // @[Mux.scala 19:72:@40604.4]
  assign inputPriorityPorts_0_5 = _T_96020[5]; // @[Mux.scala 19:72:@40606.4]
  assign inputPriorityPorts_0_6 = _T_96020[6]; // @[Mux.scala 19:72:@40608.4]
  assign inputPriorityPorts_0_7 = _T_96020[7]; // @[Mux.scala 19:72:@40610.4]
  assign inputPriorityPorts_0_8 = _T_96020[8]; // @[Mux.scala 19:72:@40612.4]
  assign inputPriorityPorts_0_9 = _T_96020[9]; // @[Mux.scala 19:72:@40614.4]
  assign inputPriorityPorts_0_10 = _T_96020[10]; // @[Mux.scala 19:72:@40616.4]
  assign inputPriorityPorts_0_11 = _T_96020[11]; // @[Mux.scala 19:72:@40618.4]
  assign inputPriorityPorts_0_12 = _T_96020[12]; // @[Mux.scala 19:72:@40620.4]
  assign inputPriorityPorts_0_13 = _T_96020[13]; // @[Mux.scala 19:72:@40622.4]
  assign inputPriorityPorts_0_14 = _T_96020[14]; // @[Mux.scala 19:72:@40624.4]
  assign inputPriorityPorts_0_15 = _T_96020[15]; // @[Mux.scala 19:72:@40626.4]
  assign _T_96222 = entriesPorts_0_15 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40680.4]
  assign _T_96223 = entriesPorts_0_14 ? 16'h4000 : _T_96222; // @[Mux.scala 31:69:@40681.4]
  assign _T_96224 = entriesPorts_0_13 ? 16'h2000 : _T_96223; // @[Mux.scala 31:69:@40682.4]
  assign _T_96225 = entriesPorts_0_12 ? 16'h1000 : _T_96224; // @[Mux.scala 31:69:@40683.4]
  assign _T_96226 = entriesPorts_0_11 ? 16'h800 : _T_96225; // @[Mux.scala 31:69:@40684.4]
  assign _T_96227 = entriesPorts_0_10 ? 16'h400 : _T_96226; // @[Mux.scala 31:69:@40685.4]
  assign _T_96228 = entriesPorts_0_9 ? 16'h200 : _T_96227; // @[Mux.scala 31:69:@40686.4]
  assign _T_96229 = entriesPorts_0_8 ? 16'h100 : _T_96228; // @[Mux.scala 31:69:@40687.4]
  assign _T_96230 = entriesPorts_0_7 ? 16'h80 : _T_96229; // @[Mux.scala 31:69:@40688.4]
  assign _T_96231 = entriesPorts_0_6 ? 16'h40 : _T_96230; // @[Mux.scala 31:69:@40689.4]
  assign _T_96232 = entriesPorts_0_5 ? 16'h20 : _T_96231; // @[Mux.scala 31:69:@40690.4]
  assign _T_96233 = entriesPorts_0_4 ? 16'h10 : _T_96232; // @[Mux.scala 31:69:@40691.4]
  assign _T_96234 = entriesPorts_0_3 ? 16'h8 : _T_96233; // @[Mux.scala 31:69:@40692.4]
  assign _T_96235 = entriesPorts_0_2 ? 16'h4 : _T_96234; // @[Mux.scala 31:69:@40693.4]
  assign _T_96236 = entriesPorts_0_1 ? 16'h2 : _T_96235; // @[Mux.scala 31:69:@40694.4]
  assign _T_96237 = entriesPorts_0_0 ? 16'h1 : _T_96236; // @[Mux.scala 31:69:@40695.4]
  assign _T_96238 = _T_96237[0]; // @[OneHot.scala 66:30:@40696.4]
  assign _T_96239 = _T_96237[1]; // @[OneHot.scala 66:30:@40697.4]
  assign _T_96240 = _T_96237[2]; // @[OneHot.scala 66:30:@40698.4]
  assign _T_96241 = _T_96237[3]; // @[OneHot.scala 66:30:@40699.4]
  assign _T_96242 = _T_96237[4]; // @[OneHot.scala 66:30:@40700.4]
  assign _T_96243 = _T_96237[5]; // @[OneHot.scala 66:30:@40701.4]
  assign _T_96244 = _T_96237[6]; // @[OneHot.scala 66:30:@40702.4]
  assign _T_96245 = _T_96237[7]; // @[OneHot.scala 66:30:@40703.4]
  assign _T_96246 = _T_96237[8]; // @[OneHot.scala 66:30:@40704.4]
  assign _T_96247 = _T_96237[9]; // @[OneHot.scala 66:30:@40705.4]
  assign _T_96248 = _T_96237[10]; // @[OneHot.scala 66:30:@40706.4]
  assign _T_96249 = _T_96237[11]; // @[OneHot.scala 66:30:@40707.4]
  assign _T_96250 = _T_96237[12]; // @[OneHot.scala 66:30:@40708.4]
  assign _T_96251 = _T_96237[13]; // @[OneHot.scala 66:30:@40709.4]
  assign _T_96252 = _T_96237[14]; // @[OneHot.scala 66:30:@40710.4]
  assign _T_96253 = _T_96237[15]; // @[OneHot.scala 66:30:@40711.4]
  assign _T_96294 = entriesPorts_0_0 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40729.4]
  assign _T_96295 = entriesPorts_0_15 ? 16'h4000 : _T_96294; // @[Mux.scala 31:69:@40730.4]
  assign _T_96296 = entriesPorts_0_14 ? 16'h2000 : _T_96295; // @[Mux.scala 31:69:@40731.4]
  assign _T_96297 = entriesPorts_0_13 ? 16'h1000 : _T_96296; // @[Mux.scala 31:69:@40732.4]
  assign _T_96298 = entriesPorts_0_12 ? 16'h800 : _T_96297; // @[Mux.scala 31:69:@40733.4]
  assign _T_96299 = entriesPorts_0_11 ? 16'h400 : _T_96298; // @[Mux.scala 31:69:@40734.4]
  assign _T_96300 = entriesPorts_0_10 ? 16'h200 : _T_96299; // @[Mux.scala 31:69:@40735.4]
  assign _T_96301 = entriesPorts_0_9 ? 16'h100 : _T_96300; // @[Mux.scala 31:69:@40736.4]
  assign _T_96302 = entriesPorts_0_8 ? 16'h80 : _T_96301; // @[Mux.scala 31:69:@40737.4]
  assign _T_96303 = entriesPorts_0_7 ? 16'h40 : _T_96302; // @[Mux.scala 31:69:@40738.4]
  assign _T_96304 = entriesPorts_0_6 ? 16'h20 : _T_96303; // @[Mux.scala 31:69:@40739.4]
  assign _T_96305 = entriesPorts_0_5 ? 16'h10 : _T_96304; // @[Mux.scala 31:69:@40740.4]
  assign _T_96306 = entriesPorts_0_4 ? 16'h8 : _T_96305; // @[Mux.scala 31:69:@40741.4]
  assign _T_96307 = entriesPorts_0_3 ? 16'h4 : _T_96306; // @[Mux.scala 31:69:@40742.4]
  assign _T_96308 = entriesPorts_0_2 ? 16'h2 : _T_96307; // @[Mux.scala 31:69:@40743.4]
  assign _T_96309 = entriesPorts_0_1 ? 16'h1 : _T_96308; // @[Mux.scala 31:69:@40744.4]
  assign _T_96310 = _T_96309[0]; // @[OneHot.scala 66:30:@40745.4]
  assign _T_96311 = _T_96309[1]; // @[OneHot.scala 66:30:@40746.4]
  assign _T_96312 = _T_96309[2]; // @[OneHot.scala 66:30:@40747.4]
  assign _T_96313 = _T_96309[3]; // @[OneHot.scala 66:30:@40748.4]
  assign _T_96314 = _T_96309[4]; // @[OneHot.scala 66:30:@40749.4]
  assign _T_96315 = _T_96309[5]; // @[OneHot.scala 66:30:@40750.4]
  assign _T_96316 = _T_96309[6]; // @[OneHot.scala 66:30:@40751.4]
  assign _T_96317 = _T_96309[7]; // @[OneHot.scala 66:30:@40752.4]
  assign _T_96318 = _T_96309[8]; // @[OneHot.scala 66:30:@40753.4]
  assign _T_96319 = _T_96309[9]; // @[OneHot.scala 66:30:@40754.4]
  assign _T_96320 = _T_96309[10]; // @[OneHot.scala 66:30:@40755.4]
  assign _T_96321 = _T_96309[11]; // @[OneHot.scala 66:30:@40756.4]
  assign _T_96322 = _T_96309[12]; // @[OneHot.scala 66:30:@40757.4]
  assign _T_96323 = _T_96309[13]; // @[OneHot.scala 66:30:@40758.4]
  assign _T_96324 = _T_96309[14]; // @[OneHot.scala 66:30:@40759.4]
  assign _T_96325 = _T_96309[15]; // @[OneHot.scala 66:30:@40760.4]
  assign _T_96366 = entriesPorts_0_1 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40778.4]
  assign _T_96367 = entriesPorts_0_0 ? 16'h4000 : _T_96366; // @[Mux.scala 31:69:@40779.4]
  assign _T_96368 = entriesPorts_0_15 ? 16'h2000 : _T_96367; // @[Mux.scala 31:69:@40780.4]
  assign _T_96369 = entriesPorts_0_14 ? 16'h1000 : _T_96368; // @[Mux.scala 31:69:@40781.4]
  assign _T_96370 = entriesPorts_0_13 ? 16'h800 : _T_96369; // @[Mux.scala 31:69:@40782.4]
  assign _T_96371 = entriesPorts_0_12 ? 16'h400 : _T_96370; // @[Mux.scala 31:69:@40783.4]
  assign _T_96372 = entriesPorts_0_11 ? 16'h200 : _T_96371; // @[Mux.scala 31:69:@40784.4]
  assign _T_96373 = entriesPorts_0_10 ? 16'h100 : _T_96372; // @[Mux.scala 31:69:@40785.4]
  assign _T_96374 = entriesPorts_0_9 ? 16'h80 : _T_96373; // @[Mux.scala 31:69:@40786.4]
  assign _T_96375 = entriesPorts_0_8 ? 16'h40 : _T_96374; // @[Mux.scala 31:69:@40787.4]
  assign _T_96376 = entriesPorts_0_7 ? 16'h20 : _T_96375; // @[Mux.scala 31:69:@40788.4]
  assign _T_96377 = entriesPorts_0_6 ? 16'h10 : _T_96376; // @[Mux.scala 31:69:@40789.4]
  assign _T_96378 = entriesPorts_0_5 ? 16'h8 : _T_96377; // @[Mux.scala 31:69:@40790.4]
  assign _T_96379 = entriesPorts_0_4 ? 16'h4 : _T_96378; // @[Mux.scala 31:69:@40791.4]
  assign _T_96380 = entriesPorts_0_3 ? 16'h2 : _T_96379; // @[Mux.scala 31:69:@40792.4]
  assign _T_96381 = entriesPorts_0_2 ? 16'h1 : _T_96380; // @[Mux.scala 31:69:@40793.4]
  assign _T_96382 = _T_96381[0]; // @[OneHot.scala 66:30:@40794.4]
  assign _T_96383 = _T_96381[1]; // @[OneHot.scala 66:30:@40795.4]
  assign _T_96384 = _T_96381[2]; // @[OneHot.scala 66:30:@40796.4]
  assign _T_96385 = _T_96381[3]; // @[OneHot.scala 66:30:@40797.4]
  assign _T_96386 = _T_96381[4]; // @[OneHot.scala 66:30:@40798.4]
  assign _T_96387 = _T_96381[5]; // @[OneHot.scala 66:30:@40799.4]
  assign _T_96388 = _T_96381[6]; // @[OneHot.scala 66:30:@40800.4]
  assign _T_96389 = _T_96381[7]; // @[OneHot.scala 66:30:@40801.4]
  assign _T_96390 = _T_96381[8]; // @[OneHot.scala 66:30:@40802.4]
  assign _T_96391 = _T_96381[9]; // @[OneHot.scala 66:30:@40803.4]
  assign _T_96392 = _T_96381[10]; // @[OneHot.scala 66:30:@40804.4]
  assign _T_96393 = _T_96381[11]; // @[OneHot.scala 66:30:@40805.4]
  assign _T_96394 = _T_96381[12]; // @[OneHot.scala 66:30:@40806.4]
  assign _T_96395 = _T_96381[13]; // @[OneHot.scala 66:30:@40807.4]
  assign _T_96396 = _T_96381[14]; // @[OneHot.scala 66:30:@40808.4]
  assign _T_96397 = _T_96381[15]; // @[OneHot.scala 66:30:@40809.4]
  assign _T_96438 = entriesPorts_0_2 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40827.4]
  assign _T_96439 = entriesPorts_0_1 ? 16'h4000 : _T_96438; // @[Mux.scala 31:69:@40828.4]
  assign _T_96440 = entriesPorts_0_0 ? 16'h2000 : _T_96439; // @[Mux.scala 31:69:@40829.4]
  assign _T_96441 = entriesPorts_0_15 ? 16'h1000 : _T_96440; // @[Mux.scala 31:69:@40830.4]
  assign _T_96442 = entriesPorts_0_14 ? 16'h800 : _T_96441; // @[Mux.scala 31:69:@40831.4]
  assign _T_96443 = entriesPorts_0_13 ? 16'h400 : _T_96442; // @[Mux.scala 31:69:@40832.4]
  assign _T_96444 = entriesPorts_0_12 ? 16'h200 : _T_96443; // @[Mux.scala 31:69:@40833.4]
  assign _T_96445 = entriesPorts_0_11 ? 16'h100 : _T_96444; // @[Mux.scala 31:69:@40834.4]
  assign _T_96446 = entriesPorts_0_10 ? 16'h80 : _T_96445; // @[Mux.scala 31:69:@40835.4]
  assign _T_96447 = entriesPorts_0_9 ? 16'h40 : _T_96446; // @[Mux.scala 31:69:@40836.4]
  assign _T_96448 = entriesPorts_0_8 ? 16'h20 : _T_96447; // @[Mux.scala 31:69:@40837.4]
  assign _T_96449 = entriesPorts_0_7 ? 16'h10 : _T_96448; // @[Mux.scala 31:69:@40838.4]
  assign _T_96450 = entriesPorts_0_6 ? 16'h8 : _T_96449; // @[Mux.scala 31:69:@40839.4]
  assign _T_96451 = entriesPorts_0_5 ? 16'h4 : _T_96450; // @[Mux.scala 31:69:@40840.4]
  assign _T_96452 = entriesPorts_0_4 ? 16'h2 : _T_96451; // @[Mux.scala 31:69:@40841.4]
  assign _T_96453 = entriesPorts_0_3 ? 16'h1 : _T_96452; // @[Mux.scala 31:69:@40842.4]
  assign _T_96454 = _T_96453[0]; // @[OneHot.scala 66:30:@40843.4]
  assign _T_96455 = _T_96453[1]; // @[OneHot.scala 66:30:@40844.4]
  assign _T_96456 = _T_96453[2]; // @[OneHot.scala 66:30:@40845.4]
  assign _T_96457 = _T_96453[3]; // @[OneHot.scala 66:30:@40846.4]
  assign _T_96458 = _T_96453[4]; // @[OneHot.scala 66:30:@40847.4]
  assign _T_96459 = _T_96453[5]; // @[OneHot.scala 66:30:@40848.4]
  assign _T_96460 = _T_96453[6]; // @[OneHot.scala 66:30:@40849.4]
  assign _T_96461 = _T_96453[7]; // @[OneHot.scala 66:30:@40850.4]
  assign _T_96462 = _T_96453[8]; // @[OneHot.scala 66:30:@40851.4]
  assign _T_96463 = _T_96453[9]; // @[OneHot.scala 66:30:@40852.4]
  assign _T_96464 = _T_96453[10]; // @[OneHot.scala 66:30:@40853.4]
  assign _T_96465 = _T_96453[11]; // @[OneHot.scala 66:30:@40854.4]
  assign _T_96466 = _T_96453[12]; // @[OneHot.scala 66:30:@40855.4]
  assign _T_96467 = _T_96453[13]; // @[OneHot.scala 66:30:@40856.4]
  assign _T_96468 = _T_96453[14]; // @[OneHot.scala 66:30:@40857.4]
  assign _T_96469 = _T_96453[15]; // @[OneHot.scala 66:30:@40858.4]
  assign _T_96510 = entriesPorts_0_3 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40876.4]
  assign _T_96511 = entriesPorts_0_2 ? 16'h4000 : _T_96510; // @[Mux.scala 31:69:@40877.4]
  assign _T_96512 = entriesPorts_0_1 ? 16'h2000 : _T_96511; // @[Mux.scala 31:69:@40878.4]
  assign _T_96513 = entriesPorts_0_0 ? 16'h1000 : _T_96512; // @[Mux.scala 31:69:@40879.4]
  assign _T_96514 = entriesPorts_0_15 ? 16'h800 : _T_96513; // @[Mux.scala 31:69:@40880.4]
  assign _T_96515 = entriesPorts_0_14 ? 16'h400 : _T_96514; // @[Mux.scala 31:69:@40881.4]
  assign _T_96516 = entriesPorts_0_13 ? 16'h200 : _T_96515; // @[Mux.scala 31:69:@40882.4]
  assign _T_96517 = entriesPorts_0_12 ? 16'h100 : _T_96516; // @[Mux.scala 31:69:@40883.4]
  assign _T_96518 = entriesPorts_0_11 ? 16'h80 : _T_96517; // @[Mux.scala 31:69:@40884.4]
  assign _T_96519 = entriesPorts_0_10 ? 16'h40 : _T_96518; // @[Mux.scala 31:69:@40885.4]
  assign _T_96520 = entriesPorts_0_9 ? 16'h20 : _T_96519; // @[Mux.scala 31:69:@40886.4]
  assign _T_96521 = entriesPorts_0_8 ? 16'h10 : _T_96520; // @[Mux.scala 31:69:@40887.4]
  assign _T_96522 = entriesPorts_0_7 ? 16'h8 : _T_96521; // @[Mux.scala 31:69:@40888.4]
  assign _T_96523 = entriesPorts_0_6 ? 16'h4 : _T_96522; // @[Mux.scala 31:69:@40889.4]
  assign _T_96524 = entriesPorts_0_5 ? 16'h2 : _T_96523; // @[Mux.scala 31:69:@40890.4]
  assign _T_96525 = entriesPorts_0_4 ? 16'h1 : _T_96524; // @[Mux.scala 31:69:@40891.4]
  assign _T_96526 = _T_96525[0]; // @[OneHot.scala 66:30:@40892.4]
  assign _T_96527 = _T_96525[1]; // @[OneHot.scala 66:30:@40893.4]
  assign _T_96528 = _T_96525[2]; // @[OneHot.scala 66:30:@40894.4]
  assign _T_96529 = _T_96525[3]; // @[OneHot.scala 66:30:@40895.4]
  assign _T_96530 = _T_96525[4]; // @[OneHot.scala 66:30:@40896.4]
  assign _T_96531 = _T_96525[5]; // @[OneHot.scala 66:30:@40897.4]
  assign _T_96532 = _T_96525[6]; // @[OneHot.scala 66:30:@40898.4]
  assign _T_96533 = _T_96525[7]; // @[OneHot.scala 66:30:@40899.4]
  assign _T_96534 = _T_96525[8]; // @[OneHot.scala 66:30:@40900.4]
  assign _T_96535 = _T_96525[9]; // @[OneHot.scala 66:30:@40901.4]
  assign _T_96536 = _T_96525[10]; // @[OneHot.scala 66:30:@40902.4]
  assign _T_96537 = _T_96525[11]; // @[OneHot.scala 66:30:@40903.4]
  assign _T_96538 = _T_96525[12]; // @[OneHot.scala 66:30:@40904.4]
  assign _T_96539 = _T_96525[13]; // @[OneHot.scala 66:30:@40905.4]
  assign _T_96540 = _T_96525[14]; // @[OneHot.scala 66:30:@40906.4]
  assign _T_96541 = _T_96525[15]; // @[OneHot.scala 66:30:@40907.4]
  assign _T_96582 = entriesPorts_0_4 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40925.4]
  assign _T_96583 = entriesPorts_0_3 ? 16'h4000 : _T_96582; // @[Mux.scala 31:69:@40926.4]
  assign _T_96584 = entriesPorts_0_2 ? 16'h2000 : _T_96583; // @[Mux.scala 31:69:@40927.4]
  assign _T_96585 = entriesPorts_0_1 ? 16'h1000 : _T_96584; // @[Mux.scala 31:69:@40928.4]
  assign _T_96586 = entriesPorts_0_0 ? 16'h800 : _T_96585; // @[Mux.scala 31:69:@40929.4]
  assign _T_96587 = entriesPorts_0_15 ? 16'h400 : _T_96586; // @[Mux.scala 31:69:@40930.4]
  assign _T_96588 = entriesPorts_0_14 ? 16'h200 : _T_96587; // @[Mux.scala 31:69:@40931.4]
  assign _T_96589 = entriesPorts_0_13 ? 16'h100 : _T_96588; // @[Mux.scala 31:69:@40932.4]
  assign _T_96590 = entriesPorts_0_12 ? 16'h80 : _T_96589; // @[Mux.scala 31:69:@40933.4]
  assign _T_96591 = entriesPorts_0_11 ? 16'h40 : _T_96590; // @[Mux.scala 31:69:@40934.4]
  assign _T_96592 = entriesPorts_0_10 ? 16'h20 : _T_96591; // @[Mux.scala 31:69:@40935.4]
  assign _T_96593 = entriesPorts_0_9 ? 16'h10 : _T_96592; // @[Mux.scala 31:69:@40936.4]
  assign _T_96594 = entriesPorts_0_8 ? 16'h8 : _T_96593; // @[Mux.scala 31:69:@40937.4]
  assign _T_96595 = entriesPorts_0_7 ? 16'h4 : _T_96594; // @[Mux.scala 31:69:@40938.4]
  assign _T_96596 = entriesPorts_0_6 ? 16'h2 : _T_96595; // @[Mux.scala 31:69:@40939.4]
  assign _T_96597 = entriesPorts_0_5 ? 16'h1 : _T_96596; // @[Mux.scala 31:69:@40940.4]
  assign _T_96598 = _T_96597[0]; // @[OneHot.scala 66:30:@40941.4]
  assign _T_96599 = _T_96597[1]; // @[OneHot.scala 66:30:@40942.4]
  assign _T_96600 = _T_96597[2]; // @[OneHot.scala 66:30:@40943.4]
  assign _T_96601 = _T_96597[3]; // @[OneHot.scala 66:30:@40944.4]
  assign _T_96602 = _T_96597[4]; // @[OneHot.scala 66:30:@40945.4]
  assign _T_96603 = _T_96597[5]; // @[OneHot.scala 66:30:@40946.4]
  assign _T_96604 = _T_96597[6]; // @[OneHot.scala 66:30:@40947.4]
  assign _T_96605 = _T_96597[7]; // @[OneHot.scala 66:30:@40948.4]
  assign _T_96606 = _T_96597[8]; // @[OneHot.scala 66:30:@40949.4]
  assign _T_96607 = _T_96597[9]; // @[OneHot.scala 66:30:@40950.4]
  assign _T_96608 = _T_96597[10]; // @[OneHot.scala 66:30:@40951.4]
  assign _T_96609 = _T_96597[11]; // @[OneHot.scala 66:30:@40952.4]
  assign _T_96610 = _T_96597[12]; // @[OneHot.scala 66:30:@40953.4]
  assign _T_96611 = _T_96597[13]; // @[OneHot.scala 66:30:@40954.4]
  assign _T_96612 = _T_96597[14]; // @[OneHot.scala 66:30:@40955.4]
  assign _T_96613 = _T_96597[15]; // @[OneHot.scala 66:30:@40956.4]
  assign _T_96654 = entriesPorts_0_5 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40974.4]
  assign _T_96655 = entriesPorts_0_4 ? 16'h4000 : _T_96654; // @[Mux.scala 31:69:@40975.4]
  assign _T_96656 = entriesPorts_0_3 ? 16'h2000 : _T_96655; // @[Mux.scala 31:69:@40976.4]
  assign _T_96657 = entriesPorts_0_2 ? 16'h1000 : _T_96656; // @[Mux.scala 31:69:@40977.4]
  assign _T_96658 = entriesPorts_0_1 ? 16'h800 : _T_96657; // @[Mux.scala 31:69:@40978.4]
  assign _T_96659 = entriesPorts_0_0 ? 16'h400 : _T_96658; // @[Mux.scala 31:69:@40979.4]
  assign _T_96660 = entriesPorts_0_15 ? 16'h200 : _T_96659; // @[Mux.scala 31:69:@40980.4]
  assign _T_96661 = entriesPorts_0_14 ? 16'h100 : _T_96660; // @[Mux.scala 31:69:@40981.4]
  assign _T_96662 = entriesPorts_0_13 ? 16'h80 : _T_96661; // @[Mux.scala 31:69:@40982.4]
  assign _T_96663 = entriesPorts_0_12 ? 16'h40 : _T_96662; // @[Mux.scala 31:69:@40983.4]
  assign _T_96664 = entriesPorts_0_11 ? 16'h20 : _T_96663; // @[Mux.scala 31:69:@40984.4]
  assign _T_96665 = entriesPorts_0_10 ? 16'h10 : _T_96664; // @[Mux.scala 31:69:@40985.4]
  assign _T_96666 = entriesPorts_0_9 ? 16'h8 : _T_96665; // @[Mux.scala 31:69:@40986.4]
  assign _T_96667 = entriesPorts_0_8 ? 16'h4 : _T_96666; // @[Mux.scala 31:69:@40987.4]
  assign _T_96668 = entriesPorts_0_7 ? 16'h2 : _T_96667; // @[Mux.scala 31:69:@40988.4]
  assign _T_96669 = entriesPorts_0_6 ? 16'h1 : _T_96668; // @[Mux.scala 31:69:@40989.4]
  assign _T_96670 = _T_96669[0]; // @[OneHot.scala 66:30:@40990.4]
  assign _T_96671 = _T_96669[1]; // @[OneHot.scala 66:30:@40991.4]
  assign _T_96672 = _T_96669[2]; // @[OneHot.scala 66:30:@40992.4]
  assign _T_96673 = _T_96669[3]; // @[OneHot.scala 66:30:@40993.4]
  assign _T_96674 = _T_96669[4]; // @[OneHot.scala 66:30:@40994.4]
  assign _T_96675 = _T_96669[5]; // @[OneHot.scala 66:30:@40995.4]
  assign _T_96676 = _T_96669[6]; // @[OneHot.scala 66:30:@40996.4]
  assign _T_96677 = _T_96669[7]; // @[OneHot.scala 66:30:@40997.4]
  assign _T_96678 = _T_96669[8]; // @[OneHot.scala 66:30:@40998.4]
  assign _T_96679 = _T_96669[9]; // @[OneHot.scala 66:30:@40999.4]
  assign _T_96680 = _T_96669[10]; // @[OneHot.scala 66:30:@41000.4]
  assign _T_96681 = _T_96669[11]; // @[OneHot.scala 66:30:@41001.4]
  assign _T_96682 = _T_96669[12]; // @[OneHot.scala 66:30:@41002.4]
  assign _T_96683 = _T_96669[13]; // @[OneHot.scala 66:30:@41003.4]
  assign _T_96684 = _T_96669[14]; // @[OneHot.scala 66:30:@41004.4]
  assign _T_96685 = _T_96669[15]; // @[OneHot.scala 66:30:@41005.4]
  assign _T_96726 = entriesPorts_0_6 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41023.4]
  assign _T_96727 = entriesPorts_0_5 ? 16'h4000 : _T_96726; // @[Mux.scala 31:69:@41024.4]
  assign _T_96728 = entriesPorts_0_4 ? 16'h2000 : _T_96727; // @[Mux.scala 31:69:@41025.4]
  assign _T_96729 = entriesPorts_0_3 ? 16'h1000 : _T_96728; // @[Mux.scala 31:69:@41026.4]
  assign _T_96730 = entriesPorts_0_2 ? 16'h800 : _T_96729; // @[Mux.scala 31:69:@41027.4]
  assign _T_96731 = entriesPorts_0_1 ? 16'h400 : _T_96730; // @[Mux.scala 31:69:@41028.4]
  assign _T_96732 = entriesPorts_0_0 ? 16'h200 : _T_96731; // @[Mux.scala 31:69:@41029.4]
  assign _T_96733 = entriesPorts_0_15 ? 16'h100 : _T_96732; // @[Mux.scala 31:69:@41030.4]
  assign _T_96734 = entriesPorts_0_14 ? 16'h80 : _T_96733; // @[Mux.scala 31:69:@41031.4]
  assign _T_96735 = entriesPorts_0_13 ? 16'h40 : _T_96734; // @[Mux.scala 31:69:@41032.4]
  assign _T_96736 = entriesPorts_0_12 ? 16'h20 : _T_96735; // @[Mux.scala 31:69:@41033.4]
  assign _T_96737 = entriesPorts_0_11 ? 16'h10 : _T_96736; // @[Mux.scala 31:69:@41034.4]
  assign _T_96738 = entriesPorts_0_10 ? 16'h8 : _T_96737; // @[Mux.scala 31:69:@41035.4]
  assign _T_96739 = entriesPorts_0_9 ? 16'h4 : _T_96738; // @[Mux.scala 31:69:@41036.4]
  assign _T_96740 = entriesPorts_0_8 ? 16'h2 : _T_96739; // @[Mux.scala 31:69:@41037.4]
  assign _T_96741 = entriesPorts_0_7 ? 16'h1 : _T_96740; // @[Mux.scala 31:69:@41038.4]
  assign _T_96742 = _T_96741[0]; // @[OneHot.scala 66:30:@41039.4]
  assign _T_96743 = _T_96741[1]; // @[OneHot.scala 66:30:@41040.4]
  assign _T_96744 = _T_96741[2]; // @[OneHot.scala 66:30:@41041.4]
  assign _T_96745 = _T_96741[3]; // @[OneHot.scala 66:30:@41042.4]
  assign _T_96746 = _T_96741[4]; // @[OneHot.scala 66:30:@41043.4]
  assign _T_96747 = _T_96741[5]; // @[OneHot.scala 66:30:@41044.4]
  assign _T_96748 = _T_96741[6]; // @[OneHot.scala 66:30:@41045.4]
  assign _T_96749 = _T_96741[7]; // @[OneHot.scala 66:30:@41046.4]
  assign _T_96750 = _T_96741[8]; // @[OneHot.scala 66:30:@41047.4]
  assign _T_96751 = _T_96741[9]; // @[OneHot.scala 66:30:@41048.4]
  assign _T_96752 = _T_96741[10]; // @[OneHot.scala 66:30:@41049.4]
  assign _T_96753 = _T_96741[11]; // @[OneHot.scala 66:30:@41050.4]
  assign _T_96754 = _T_96741[12]; // @[OneHot.scala 66:30:@41051.4]
  assign _T_96755 = _T_96741[13]; // @[OneHot.scala 66:30:@41052.4]
  assign _T_96756 = _T_96741[14]; // @[OneHot.scala 66:30:@41053.4]
  assign _T_96757 = _T_96741[15]; // @[OneHot.scala 66:30:@41054.4]
  assign _T_96798 = entriesPorts_0_7 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41072.4]
  assign _T_96799 = entriesPorts_0_6 ? 16'h4000 : _T_96798; // @[Mux.scala 31:69:@41073.4]
  assign _T_96800 = entriesPorts_0_5 ? 16'h2000 : _T_96799; // @[Mux.scala 31:69:@41074.4]
  assign _T_96801 = entriesPorts_0_4 ? 16'h1000 : _T_96800; // @[Mux.scala 31:69:@41075.4]
  assign _T_96802 = entriesPorts_0_3 ? 16'h800 : _T_96801; // @[Mux.scala 31:69:@41076.4]
  assign _T_96803 = entriesPorts_0_2 ? 16'h400 : _T_96802; // @[Mux.scala 31:69:@41077.4]
  assign _T_96804 = entriesPorts_0_1 ? 16'h200 : _T_96803; // @[Mux.scala 31:69:@41078.4]
  assign _T_96805 = entriesPorts_0_0 ? 16'h100 : _T_96804; // @[Mux.scala 31:69:@41079.4]
  assign _T_96806 = entriesPorts_0_15 ? 16'h80 : _T_96805; // @[Mux.scala 31:69:@41080.4]
  assign _T_96807 = entriesPorts_0_14 ? 16'h40 : _T_96806; // @[Mux.scala 31:69:@41081.4]
  assign _T_96808 = entriesPorts_0_13 ? 16'h20 : _T_96807; // @[Mux.scala 31:69:@41082.4]
  assign _T_96809 = entriesPorts_0_12 ? 16'h10 : _T_96808; // @[Mux.scala 31:69:@41083.4]
  assign _T_96810 = entriesPorts_0_11 ? 16'h8 : _T_96809; // @[Mux.scala 31:69:@41084.4]
  assign _T_96811 = entriesPorts_0_10 ? 16'h4 : _T_96810; // @[Mux.scala 31:69:@41085.4]
  assign _T_96812 = entriesPorts_0_9 ? 16'h2 : _T_96811; // @[Mux.scala 31:69:@41086.4]
  assign _T_96813 = entriesPorts_0_8 ? 16'h1 : _T_96812; // @[Mux.scala 31:69:@41087.4]
  assign _T_96814 = _T_96813[0]; // @[OneHot.scala 66:30:@41088.4]
  assign _T_96815 = _T_96813[1]; // @[OneHot.scala 66:30:@41089.4]
  assign _T_96816 = _T_96813[2]; // @[OneHot.scala 66:30:@41090.4]
  assign _T_96817 = _T_96813[3]; // @[OneHot.scala 66:30:@41091.4]
  assign _T_96818 = _T_96813[4]; // @[OneHot.scala 66:30:@41092.4]
  assign _T_96819 = _T_96813[5]; // @[OneHot.scala 66:30:@41093.4]
  assign _T_96820 = _T_96813[6]; // @[OneHot.scala 66:30:@41094.4]
  assign _T_96821 = _T_96813[7]; // @[OneHot.scala 66:30:@41095.4]
  assign _T_96822 = _T_96813[8]; // @[OneHot.scala 66:30:@41096.4]
  assign _T_96823 = _T_96813[9]; // @[OneHot.scala 66:30:@41097.4]
  assign _T_96824 = _T_96813[10]; // @[OneHot.scala 66:30:@41098.4]
  assign _T_96825 = _T_96813[11]; // @[OneHot.scala 66:30:@41099.4]
  assign _T_96826 = _T_96813[12]; // @[OneHot.scala 66:30:@41100.4]
  assign _T_96827 = _T_96813[13]; // @[OneHot.scala 66:30:@41101.4]
  assign _T_96828 = _T_96813[14]; // @[OneHot.scala 66:30:@41102.4]
  assign _T_96829 = _T_96813[15]; // @[OneHot.scala 66:30:@41103.4]
  assign _T_96870 = entriesPorts_0_8 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41121.4]
  assign _T_96871 = entriesPorts_0_7 ? 16'h4000 : _T_96870; // @[Mux.scala 31:69:@41122.4]
  assign _T_96872 = entriesPorts_0_6 ? 16'h2000 : _T_96871; // @[Mux.scala 31:69:@41123.4]
  assign _T_96873 = entriesPorts_0_5 ? 16'h1000 : _T_96872; // @[Mux.scala 31:69:@41124.4]
  assign _T_96874 = entriesPorts_0_4 ? 16'h800 : _T_96873; // @[Mux.scala 31:69:@41125.4]
  assign _T_96875 = entriesPorts_0_3 ? 16'h400 : _T_96874; // @[Mux.scala 31:69:@41126.4]
  assign _T_96876 = entriesPorts_0_2 ? 16'h200 : _T_96875; // @[Mux.scala 31:69:@41127.4]
  assign _T_96877 = entriesPorts_0_1 ? 16'h100 : _T_96876; // @[Mux.scala 31:69:@41128.4]
  assign _T_96878 = entriesPorts_0_0 ? 16'h80 : _T_96877; // @[Mux.scala 31:69:@41129.4]
  assign _T_96879 = entriesPorts_0_15 ? 16'h40 : _T_96878; // @[Mux.scala 31:69:@41130.4]
  assign _T_96880 = entriesPorts_0_14 ? 16'h20 : _T_96879; // @[Mux.scala 31:69:@41131.4]
  assign _T_96881 = entriesPorts_0_13 ? 16'h10 : _T_96880; // @[Mux.scala 31:69:@41132.4]
  assign _T_96882 = entriesPorts_0_12 ? 16'h8 : _T_96881; // @[Mux.scala 31:69:@41133.4]
  assign _T_96883 = entriesPorts_0_11 ? 16'h4 : _T_96882; // @[Mux.scala 31:69:@41134.4]
  assign _T_96884 = entriesPorts_0_10 ? 16'h2 : _T_96883; // @[Mux.scala 31:69:@41135.4]
  assign _T_96885 = entriesPorts_0_9 ? 16'h1 : _T_96884; // @[Mux.scala 31:69:@41136.4]
  assign _T_96886 = _T_96885[0]; // @[OneHot.scala 66:30:@41137.4]
  assign _T_96887 = _T_96885[1]; // @[OneHot.scala 66:30:@41138.4]
  assign _T_96888 = _T_96885[2]; // @[OneHot.scala 66:30:@41139.4]
  assign _T_96889 = _T_96885[3]; // @[OneHot.scala 66:30:@41140.4]
  assign _T_96890 = _T_96885[4]; // @[OneHot.scala 66:30:@41141.4]
  assign _T_96891 = _T_96885[5]; // @[OneHot.scala 66:30:@41142.4]
  assign _T_96892 = _T_96885[6]; // @[OneHot.scala 66:30:@41143.4]
  assign _T_96893 = _T_96885[7]; // @[OneHot.scala 66:30:@41144.4]
  assign _T_96894 = _T_96885[8]; // @[OneHot.scala 66:30:@41145.4]
  assign _T_96895 = _T_96885[9]; // @[OneHot.scala 66:30:@41146.4]
  assign _T_96896 = _T_96885[10]; // @[OneHot.scala 66:30:@41147.4]
  assign _T_96897 = _T_96885[11]; // @[OneHot.scala 66:30:@41148.4]
  assign _T_96898 = _T_96885[12]; // @[OneHot.scala 66:30:@41149.4]
  assign _T_96899 = _T_96885[13]; // @[OneHot.scala 66:30:@41150.4]
  assign _T_96900 = _T_96885[14]; // @[OneHot.scala 66:30:@41151.4]
  assign _T_96901 = _T_96885[15]; // @[OneHot.scala 66:30:@41152.4]
  assign _T_96942 = entriesPorts_0_9 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41170.4]
  assign _T_96943 = entriesPorts_0_8 ? 16'h4000 : _T_96942; // @[Mux.scala 31:69:@41171.4]
  assign _T_96944 = entriesPorts_0_7 ? 16'h2000 : _T_96943; // @[Mux.scala 31:69:@41172.4]
  assign _T_96945 = entriesPorts_0_6 ? 16'h1000 : _T_96944; // @[Mux.scala 31:69:@41173.4]
  assign _T_96946 = entriesPorts_0_5 ? 16'h800 : _T_96945; // @[Mux.scala 31:69:@41174.4]
  assign _T_96947 = entriesPorts_0_4 ? 16'h400 : _T_96946; // @[Mux.scala 31:69:@41175.4]
  assign _T_96948 = entriesPorts_0_3 ? 16'h200 : _T_96947; // @[Mux.scala 31:69:@41176.4]
  assign _T_96949 = entriesPorts_0_2 ? 16'h100 : _T_96948; // @[Mux.scala 31:69:@41177.4]
  assign _T_96950 = entriesPorts_0_1 ? 16'h80 : _T_96949; // @[Mux.scala 31:69:@41178.4]
  assign _T_96951 = entriesPorts_0_0 ? 16'h40 : _T_96950; // @[Mux.scala 31:69:@41179.4]
  assign _T_96952 = entriesPorts_0_15 ? 16'h20 : _T_96951; // @[Mux.scala 31:69:@41180.4]
  assign _T_96953 = entriesPorts_0_14 ? 16'h10 : _T_96952; // @[Mux.scala 31:69:@41181.4]
  assign _T_96954 = entriesPorts_0_13 ? 16'h8 : _T_96953; // @[Mux.scala 31:69:@41182.4]
  assign _T_96955 = entriesPorts_0_12 ? 16'h4 : _T_96954; // @[Mux.scala 31:69:@41183.4]
  assign _T_96956 = entriesPorts_0_11 ? 16'h2 : _T_96955; // @[Mux.scala 31:69:@41184.4]
  assign _T_96957 = entriesPorts_0_10 ? 16'h1 : _T_96956; // @[Mux.scala 31:69:@41185.4]
  assign _T_96958 = _T_96957[0]; // @[OneHot.scala 66:30:@41186.4]
  assign _T_96959 = _T_96957[1]; // @[OneHot.scala 66:30:@41187.4]
  assign _T_96960 = _T_96957[2]; // @[OneHot.scala 66:30:@41188.4]
  assign _T_96961 = _T_96957[3]; // @[OneHot.scala 66:30:@41189.4]
  assign _T_96962 = _T_96957[4]; // @[OneHot.scala 66:30:@41190.4]
  assign _T_96963 = _T_96957[5]; // @[OneHot.scala 66:30:@41191.4]
  assign _T_96964 = _T_96957[6]; // @[OneHot.scala 66:30:@41192.4]
  assign _T_96965 = _T_96957[7]; // @[OneHot.scala 66:30:@41193.4]
  assign _T_96966 = _T_96957[8]; // @[OneHot.scala 66:30:@41194.4]
  assign _T_96967 = _T_96957[9]; // @[OneHot.scala 66:30:@41195.4]
  assign _T_96968 = _T_96957[10]; // @[OneHot.scala 66:30:@41196.4]
  assign _T_96969 = _T_96957[11]; // @[OneHot.scala 66:30:@41197.4]
  assign _T_96970 = _T_96957[12]; // @[OneHot.scala 66:30:@41198.4]
  assign _T_96971 = _T_96957[13]; // @[OneHot.scala 66:30:@41199.4]
  assign _T_96972 = _T_96957[14]; // @[OneHot.scala 66:30:@41200.4]
  assign _T_96973 = _T_96957[15]; // @[OneHot.scala 66:30:@41201.4]
  assign _T_97014 = entriesPorts_0_10 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41219.4]
  assign _T_97015 = entriesPorts_0_9 ? 16'h4000 : _T_97014; // @[Mux.scala 31:69:@41220.4]
  assign _T_97016 = entriesPorts_0_8 ? 16'h2000 : _T_97015; // @[Mux.scala 31:69:@41221.4]
  assign _T_97017 = entriesPorts_0_7 ? 16'h1000 : _T_97016; // @[Mux.scala 31:69:@41222.4]
  assign _T_97018 = entriesPorts_0_6 ? 16'h800 : _T_97017; // @[Mux.scala 31:69:@41223.4]
  assign _T_97019 = entriesPorts_0_5 ? 16'h400 : _T_97018; // @[Mux.scala 31:69:@41224.4]
  assign _T_97020 = entriesPorts_0_4 ? 16'h200 : _T_97019; // @[Mux.scala 31:69:@41225.4]
  assign _T_97021 = entriesPorts_0_3 ? 16'h100 : _T_97020; // @[Mux.scala 31:69:@41226.4]
  assign _T_97022 = entriesPorts_0_2 ? 16'h80 : _T_97021; // @[Mux.scala 31:69:@41227.4]
  assign _T_97023 = entriesPorts_0_1 ? 16'h40 : _T_97022; // @[Mux.scala 31:69:@41228.4]
  assign _T_97024 = entriesPorts_0_0 ? 16'h20 : _T_97023; // @[Mux.scala 31:69:@41229.4]
  assign _T_97025 = entriesPorts_0_15 ? 16'h10 : _T_97024; // @[Mux.scala 31:69:@41230.4]
  assign _T_97026 = entriesPorts_0_14 ? 16'h8 : _T_97025; // @[Mux.scala 31:69:@41231.4]
  assign _T_97027 = entriesPorts_0_13 ? 16'h4 : _T_97026; // @[Mux.scala 31:69:@41232.4]
  assign _T_97028 = entriesPorts_0_12 ? 16'h2 : _T_97027; // @[Mux.scala 31:69:@41233.4]
  assign _T_97029 = entriesPorts_0_11 ? 16'h1 : _T_97028; // @[Mux.scala 31:69:@41234.4]
  assign _T_97030 = _T_97029[0]; // @[OneHot.scala 66:30:@41235.4]
  assign _T_97031 = _T_97029[1]; // @[OneHot.scala 66:30:@41236.4]
  assign _T_97032 = _T_97029[2]; // @[OneHot.scala 66:30:@41237.4]
  assign _T_97033 = _T_97029[3]; // @[OneHot.scala 66:30:@41238.4]
  assign _T_97034 = _T_97029[4]; // @[OneHot.scala 66:30:@41239.4]
  assign _T_97035 = _T_97029[5]; // @[OneHot.scala 66:30:@41240.4]
  assign _T_97036 = _T_97029[6]; // @[OneHot.scala 66:30:@41241.4]
  assign _T_97037 = _T_97029[7]; // @[OneHot.scala 66:30:@41242.4]
  assign _T_97038 = _T_97029[8]; // @[OneHot.scala 66:30:@41243.4]
  assign _T_97039 = _T_97029[9]; // @[OneHot.scala 66:30:@41244.4]
  assign _T_97040 = _T_97029[10]; // @[OneHot.scala 66:30:@41245.4]
  assign _T_97041 = _T_97029[11]; // @[OneHot.scala 66:30:@41246.4]
  assign _T_97042 = _T_97029[12]; // @[OneHot.scala 66:30:@41247.4]
  assign _T_97043 = _T_97029[13]; // @[OneHot.scala 66:30:@41248.4]
  assign _T_97044 = _T_97029[14]; // @[OneHot.scala 66:30:@41249.4]
  assign _T_97045 = _T_97029[15]; // @[OneHot.scala 66:30:@41250.4]
  assign _T_97086 = entriesPorts_0_11 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41268.4]
  assign _T_97087 = entriesPorts_0_10 ? 16'h4000 : _T_97086; // @[Mux.scala 31:69:@41269.4]
  assign _T_97088 = entriesPorts_0_9 ? 16'h2000 : _T_97087; // @[Mux.scala 31:69:@41270.4]
  assign _T_97089 = entriesPorts_0_8 ? 16'h1000 : _T_97088; // @[Mux.scala 31:69:@41271.4]
  assign _T_97090 = entriesPorts_0_7 ? 16'h800 : _T_97089; // @[Mux.scala 31:69:@41272.4]
  assign _T_97091 = entriesPorts_0_6 ? 16'h400 : _T_97090; // @[Mux.scala 31:69:@41273.4]
  assign _T_97092 = entriesPorts_0_5 ? 16'h200 : _T_97091; // @[Mux.scala 31:69:@41274.4]
  assign _T_97093 = entriesPorts_0_4 ? 16'h100 : _T_97092; // @[Mux.scala 31:69:@41275.4]
  assign _T_97094 = entriesPorts_0_3 ? 16'h80 : _T_97093; // @[Mux.scala 31:69:@41276.4]
  assign _T_97095 = entriesPorts_0_2 ? 16'h40 : _T_97094; // @[Mux.scala 31:69:@41277.4]
  assign _T_97096 = entriesPorts_0_1 ? 16'h20 : _T_97095; // @[Mux.scala 31:69:@41278.4]
  assign _T_97097 = entriesPorts_0_0 ? 16'h10 : _T_97096; // @[Mux.scala 31:69:@41279.4]
  assign _T_97098 = entriesPorts_0_15 ? 16'h8 : _T_97097; // @[Mux.scala 31:69:@41280.4]
  assign _T_97099 = entriesPorts_0_14 ? 16'h4 : _T_97098; // @[Mux.scala 31:69:@41281.4]
  assign _T_97100 = entriesPorts_0_13 ? 16'h2 : _T_97099; // @[Mux.scala 31:69:@41282.4]
  assign _T_97101 = entriesPorts_0_12 ? 16'h1 : _T_97100; // @[Mux.scala 31:69:@41283.4]
  assign _T_97102 = _T_97101[0]; // @[OneHot.scala 66:30:@41284.4]
  assign _T_97103 = _T_97101[1]; // @[OneHot.scala 66:30:@41285.4]
  assign _T_97104 = _T_97101[2]; // @[OneHot.scala 66:30:@41286.4]
  assign _T_97105 = _T_97101[3]; // @[OneHot.scala 66:30:@41287.4]
  assign _T_97106 = _T_97101[4]; // @[OneHot.scala 66:30:@41288.4]
  assign _T_97107 = _T_97101[5]; // @[OneHot.scala 66:30:@41289.4]
  assign _T_97108 = _T_97101[6]; // @[OneHot.scala 66:30:@41290.4]
  assign _T_97109 = _T_97101[7]; // @[OneHot.scala 66:30:@41291.4]
  assign _T_97110 = _T_97101[8]; // @[OneHot.scala 66:30:@41292.4]
  assign _T_97111 = _T_97101[9]; // @[OneHot.scala 66:30:@41293.4]
  assign _T_97112 = _T_97101[10]; // @[OneHot.scala 66:30:@41294.4]
  assign _T_97113 = _T_97101[11]; // @[OneHot.scala 66:30:@41295.4]
  assign _T_97114 = _T_97101[12]; // @[OneHot.scala 66:30:@41296.4]
  assign _T_97115 = _T_97101[13]; // @[OneHot.scala 66:30:@41297.4]
  assign _T_97116 = _T_97101[14]; // @[OneHot.scala 66:30:@41298.4]
  assign _T_97117 = _T_97101[15]; // @[OneHot.scala 66:30:@41299.4]
  assign _T_97158 = entriesPorts_0_12 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41317.4]
  assign _T_97159 = entriesPorts_0_11 ? 16'h4000 : _T_97158; // @[Mux.scala 31:69:@41318.4]
  assign _T_97160 = entriesPorts_0_10 ? 16'h2000 : _T_97159; // @[Mux.scala 31:69:@41319.4]
  assign _T_97161 = entriesPorts_0_9 ? 16'h1000 : _T_97160; // @[Mux.scala 31:69:@41320.4]
  assign _T_97162 = entriesPorts_0_8 ? 16'h800 : _T_97161; // @[Mux.scala 31:69:@41321.4]
  assign _T_97163 = entriesPorts_0_7 ? 16'h400 : _T_97162; // @[Mux.scala 31:69:@41322.4]
  assign _T_97164 = entriesPorts_0_6 ? 16'h200 : _T_97163; // @[Mux.scala 31:69:@41323.4]
  assign _T_97165 = entriesPorts_0_5 ? 16'h100 : _T_97164; // @[Mux.scala 31:69:@41324.4]
  assign _T_97166 = entriesPorts_0_4 ? 16'h80 : _T_97165; // @[Mux.scala 31:69:@41325.4]
  assign _T_97167 = entriesPorts_0_3 ? 16'h40 : _T_97166; // @[Mux.scala 31:69:@41326.4]
  assign _T_97168 = entriesPorts_0_2 ? 16'h20 : _T_97167; // @[Mux.scala 31:69:@41327.4]
  assign _T_97169 = entriesPorts_0_1 ? 16'h10 : _T_97168; // @[Mux.scala 31:69:@41328.4]
  assign _T_97170 = entriesPorts_0_0 ? 16'h8 : _T_97169; // @[Mux.scala 31:69:@41329.4]
  assign _T_97171 = entriesPorts_0_15 ? 16'h4 : _T_97170; // @[Mux.scala 31:69:@41330.4]
  assign _T_97172 = entriesPorts_0_14 ? 16'h2 : _T_97171; // @[Mux.scala 31:69:@41331.4]
  assign _T_97173 = entriesPorts_0_13 ? 16'h1 : _T_97172; // @[Mux.scala 31:69:@41332.4]
  assign _T_97174 = _T_97173[0]; // @[OneHot.scala 66:30:@41333.4]
  assign _T_97175 = _T_97173[1]; // @[OneHot.scala 66:30:@41334.4]
  assign _T_97176 = _T_97173[2]; // @[OneHot.scala 66:30:@41335.4]
  assign _T_97177 = _T_97173[3]; // @[OneHot.scala 66:30:@41336.4]
  assign _T_97178 = _T_97173[4]; // @[OneHot.scala 66:30:@41337.4]
  assign _T_97179 = _T_97173[5]; // @[OneHot.scala 66:30:@41338.4]
  assign _T_97180 = _T_97173[6]; // @[OneHot.scala 66:30:@41339.4]
  assign _T_97181 = _T_97173[7]; // @[OneHot.scala 66:30:@41340.4]
  assign _T_97182 = _T_97173[8]; // @[OneHot.scala 66:30:@41341.4]
  assign _T_97183 = _T_97173[9]; // @[OneHot.scala 66:30:@41342.4]
  assign _T_97184 = _T_97173[10]; // @[OneHot.scala 66:30:@41343.4]
  assign _T_97185 = _T_97173[11]; // @[OneHot.scala 66:30:@41344.4]
  assign _T_97186 = _T_97173[12]; // @[OneHot.scala 66:30:@41345.4]
  assign _T_97187 = _T_97173[13]; // @[OneHot.scala 66:30:@41346.4]
  assign _T_97188 = _T_97173[14]; // @[OneHot.scala 66:30:@41347.4]
  assign _T_97189 = _T_97173[15]; // @[OneHot.scala 66:30:@41348.4]
  assign _T_97230 = entriesPorts_0_13 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41366.4]
  assign _T_97231 = entriesPorts_0_12 ? 16'h4000 : _T_97230; // @[Mux.scala 31:69:@41367.4]
  assign _T_97232 = entriesPorts_0_11 ? 16'h2000 : _T_97231; // @[Mux.scala 31:69:@41368.4]
  assign _T_97233 = entriesPorts_0_10 ? 16'h1000 : _T_97232; // @[Mux.scala 31:69:@41369.4]
  assign _T_97234 = entriesPorts_0_9 ? 16'h800 : _T_97233; // @[Mux.scala 31:69:@41370.4]
  assign _T_97235 = entriesPorts_0_8 ? 16'h400 : _T_97234; // @[Mux.scala 31:69:@41371.4]
  assign _T_97236 = entriesPorts_0_7 ? 16'h200 : _T_97235; // @[Mux.scala 31:69:@41372.4]
  assign _T_97237 = entriesPorts_0_6 ? 16'h100 : _T_97236; // @[Mux.scala 31:69:@41373.4]
  assign _T_97238 = entriesPorts_0_5 ? 16'h80 : _T_97237; // @[Mux.scala 31:69:@41374.4]
  assign _T_97239 = entriesPorts_0_4 ? 16'h40 : _T_97238; // @[Mux.scala 31:69:@41375.4]
  assign _T_97240 = entriesPorts_0_3 ? 16'h20 : _T_97239; // @[Mux.scala 31:69:@41376.4]
  assign _T_97241 = entriesPorts_0_2 ? 16'h10 : _T_97240; // @[Mux.scala 31:69:@41377.4]
  assign _T_97242 = entriesPorts_0_1 ? 16'h8 : _T_97241; // @[Mux.scala 31:69:@41378.4]
  assign _T_97243 = entriesPorts_0_0 ? 16'h4 : _T_97242; // @[Mux.scala 31:69:@41379.4]
  assign _T_97244 = entriesPorts_0_15 ? 16'h2 : _T_97243; // @[Mux.scala 31:69:@41380.4]
  assign _T_97245 = entriesPorts_0_14 ? 16'h1 : _T_97244; // @[Mux.scala 31:69:@41381.4]
  assign _T_97246 = _T_97245[0]; // @[OneHot.scala 66:30:@41382.4]
  assign _T_97247 = _T_97245[1]; // @[OneHot.scala 66:30:@41383.4]
  assign _T_97248 = _T_97245[2]; // @[OneHot.scala 66:30:@41384.4]
  assign _T_97249 = _T_97245[3]; // @[OneHot.scala 66:30:@41385.4]
  assign _T_97250 = _T_97245[4]; // @[OneHot.scala 66:30:@41386.4]
  assign _T_97251 = _T_97245[5]; // @[OneHot.scala 66:30:@41387.4]
  assign _T_97252 = _T_97245[6]; // @[OneHot.scala 66:30:@41388.4]
  assign _T_97253 = _T_97245[7]; // @[OneHot.scala 66:30:@41389.4]
  assign _T_97254 = _T_97245[8]; // @[OneHot.scala 66:30:@41390.4]
  assign _T_97255 = _T_97245[9]; // @[OneHot.scala 66:30:@41391.4]
  assign _T_97256 = _T_97245[10]; // @[OneHot.scala 66:30:@41392.4]
  assign _T_97257 = _T_97245[11]; // @[OneHot.scala 66:30:@41393.4]
  assign _T_97258 = _T_97245[12]; // @[OneHot.scala 66:30:@41394.4]
  assign _T_97259 = _T_97245[13]; // @[OneHot.scala 66:30:@41395.4]
  assign _T_97260 = _T_97245[14]; // @[OneHot.scala 66:30:@41396.4]
  assign _T_97261 = _T_97245[15]; // @[OneHot.scala 66:30:@41397.4]
  assign _T_97302 = entriesPorts_0_14 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41415.4]
  assign _T_97303 = entriesPorts_0_13 ? 16'h4000 : _T_97302; // @[Mux.scala 31:69:@41416.4]
  assign _T_97304 = entriesPorts_0_12 ? 16'h2000 : _T_97303; // @[Mux.scala 31:69:@41417.4]
  assign _T_97305 = entriesPorts_0_11 ? 16'h1000 : _T_97304; // @[Mux.scala 31:69:@41418.4]
  assign _T_97306 = entriesPorts_0_10 ? 16'h800 : _T_97305; // @[Mux.scala 31:69:@41419.4]
  assign _T_97307 = entriesPorts_0_9 ? 16'h400 : _T_97306; // @[Mux.scala 31:69:@41420.4]
  assign _T_97308 = entriesPorts_0_8 ? 16'h200 : _T_97307; // @[Mux.scala 31:69:@41421.4]
  assign _T_97309 = entriesPorts_0_7 ? 16'h100 : _T_97308; // @[Mux.scala 31:69:@41422.4]
  assign _T_97310 = entriesPorts_0_6 ? 16'h80 : _T_97309; // @[Mux.scala 31:69:@41423.4]
  assign _T_97311 = entriesPorts_0_5 ? 16'h40 : _T_97310; // @[Mux.scala 31:69:@41424.4]
  assign _T_97312 = entriesPorts_0_4 ? 16'h20 : _T_97311; // @[Mux.scala 31:69:@41425.4]
  assign _T_97313 = entriesPorts_0_3 ? 16'h10 : _T_97312; // @[Mux.scala 31:69:@41426.4]
  assign _T_97314 = entriesPorts_0_2 ? 16'h8 : _T_97313; // @[Mux.scala 31:69:@41427.4]
  assign _T_97315 = entriesPorts_0_1 ? 16'h4 : _T_97314; // @[Mux.scala 31:69:@41428.4]
  assign _T_97316 = entriesPorts_0_0 ? 16'h2 : _T_97315; // @[Mux.scala 31:69:@41429.4]
  assign _T_97317 = entriesPorts_0_15 ? 16'h1 : _T_97316; // @[Mux.scala 31:69:@41430.4]
  assign _T_97318 = _T_97317[0]; // @[OneHot.scala 66:30:@41431.4]
  assign _T_97319 = _T_97317[1]; // @[OneHot.scala 66:30:@41432.4]
  assign _T_97320 = _T_97317[2]; // @[OneHot.scala 66:30:@41433.4]
  assign _T_97321 = _T_97317[3]; // @[OneHot.scala 66:30:@41434.4]
  assign _T_97322 = _T_97317[4]; // @[OneHot.scala 66:30:@41435.4]
  assign _T_97323 = _T_97317[5]; // @[OneHot.scala 66:30:@41436.4]
  assign _T_97324 = _T_97317[6]; // @[OneHot.scala 66:30:@41437.4]
  assign _T_97325 = _T_97317[7]; // @[OneHot.scala 66:30:@41438.4]
  assign _T_97326 = _T_97317[8]; // @[OneHot.scala 66:30:@41439.4]
  assign _T_97327 = _T_97317[9]; // @[OneHot.scala 66:30:@41440.4]
  assign _T_97328 = _T_97317[10]; // @[OneHot.scala 66:30:@41441.4]
  assign _T_97329 = _T_97317[11]; // @[OneHot.scala 66:30:@41442.4]
  assign _T_97330 = _T_97317[12]; // @[OneHot.scala 66:30:@41443.4]
  assign _T_97331 = _T_97317[13]; // @[OneHot.scala 66:30:@41444.4]
  assign _T_97332 = _T_97317[14]; // @[OneHot.scala 66:30:@41445.4]
  assign _T_97333 = _T_97317[15]; // @[OneHot.scala 66:30:@41446.4]
  assign _T_97398 = {_T_96245,_T_96244,_T_96243,_T_96242,_T_96241,_T_96240,_T_96239,_T_96238}; // @[Mux.scala 19:72:@41470.4]
  assign _T_97406 = {_T_96253,_T_96252,_T_96251,_T_96250,_T_96249,_T_96248,_T_96247,_T_96246,_T_97398}; // @[Mux.scala 19:72:@41478.4]
  assign _T_97408 = _T_90408 ? _T_97406 : 16'h0; // @[Mux.scala 19:72:@41479.4]
  assign _T_97415 = {_T_96316,_T_96315,_T_96314,_T_96313,_T_96312,_T_96311,_T_96310,_T_96325}; // @[Mux.scala 19:72:@41486.4]
  assign _T_97423 = {_T_96324,_T_96323,_T_96322,_T_96321,_T_96320,_T_96319,_T_96318,_T_96317,_T_97415}; // @[Mux.scala 19:72:@41494.4]
  assign _T_97425 = _T_90409 ? _T_97423 : 16'h0; // @[Mux.scala 19:72:@41495.4]
  assign _T_97432 = {_T_96387,_T_96386,_T_96385,_T_96384,_T_96383,_T_96382,_T_96397,_T_96396}; // @[Mux.scala 19:72:@41502.4]
  assign _T_97440 = {_T_96395,_T_96394,_T_96393,_T_96392,_T_96391,_T_96390,_T_96389,_T_96388,_T_97432}; // @[Mux.scala 19:72:@41510.4]
  assign _T_97442 = _T_90410 ? _T_97440 : 16'h0; // @[Mux.scala 19:72:@41511.4]
  assign _T_97449 = {_T_96458,_T_96457,_T_96456,_T_96455,_T_96454,_T_96469,_T_96468,_T_96467}; // @[Mux.scala 19:72:@41518.4]
  assign _T_97457 = {_T_96466,_T_96465,_T_96464,_T_96463,_T_96462,_T_96461,_T_96460,_T_96459,_T_97449}; // @[Mux.scala 19:72:@41526.4]
  assign _T_97459 = _T_90411 ? _T_97457 : 16'h0; // @[Mux.scala 19:72:@41527.4]
  assign _T_97466 = {_T_96529,_T_96528,_T_96527,_T_96526,_T_96541,_T_96540,_T_96539,_T_96538}; // @[Mux.scala 19:72:@41534.4]
  assign _T_97474 = {_T_96537,_T_96536,_T_96535,_T_96534,_T_96533,_T_96532,_T_96531,_T_96530,_T_97466}; // @[Mux.scala 19:72:@41542.4]
  assign _T_97476 = _T_90412 ? _T_97474 : 16'h0; // @[Mux.scala 19:72:@41543.4]
  assign _T_97483 = {_T_96600,_T_96599,_T_96598,_T_96613,_T_96612,_T_96611,_T_96610,_T_96609}; // @[Mux.scala 19:72:@41550.4]
  assign _T_97491 = {_T_96608,_T_96607,_T_96606,_T_96605,_T_96604,_T_96603,_T_96602,_T_96601,_T_97483}; // @[Mux.scala 19:72:@41558.4]
  assign _T_97493 = _T_90413 ? _T_97491 : 16'h0; // @[Mux.scala 19:72:@41559.4]
  assign _T_97500 = {_T_96671,_T_96670,_T_96685,_T_96684,_T_96683,_T_96682,_T_96681,_T_96680}; // @[Mux.scala 19:72:@41566.4]
  assign _T_97508 = {_T_96679,_T_96678,_T_96677,_T_96676,_T_96675,_T_96674,_T_96673,_T_96672,_T_97500}; // @[Mux.scala 19:72:@41574.4]
  assign _T_97510 = _T_90414 ? _T_97508 : 16'h0; // @[Mux.scala 19:72:@41575.4]
  assign _T_97517 = {_T_96742,_T_96757,_T_96756,_T_96755,_T_96754,_T_96753,_T_96752,_T_96751}; // @[Mux.scala 19:72:@41582.4]
  assign _T_97525 = {_T_96750,_T_96749,_T_96748,_T_96747,_T_96746,_T_96745,_T_96744,_T_96743,_T_97517}; // @[Mux.scala 19:72:@41590.4]
  assign _T_97527 = _T_90415 ? _T_97525 : 16'h0; // @[Mux.scala 19:72:@41591.4]
  assign _T_97534 = {_T_96829,_T_96828,_T_96827,_T_96826,_T_96825,_T_96824,_T_96823,_T_96822}; // @[Mux.scala 19:72:@41598.4]
  assign _T_97542 = {_T_96821,_T_96820,_T_96819,_T_96818,_T_96817,_T_96816,_T_96815,_T_96814,_T_97534}; // @[Mux.scala 19:72:@41606.4]
  assign _T_97544 = _T_90416 ? _T_97542 : 16'h0; // @[Mux.scala 19:72:@41607.4]
  assign _T_97551 = {_T_96900,_T_96899,_T_96898,_T_96897,_T_96896,_T_96895,_T_96894,_T_96893}; // @[Mux.scala 19:72:@41614.4]
  assign _T_97559 = {_T_96892,_T_96891,_T_96890,_T_96889,_T_96888,_T_96887,_T_96886,_T_96901,_T_97551}; // @[Mux.scala 19:72:@41622.4]
  assign _T_97561 = _T_90417 ? _T_97559 : 16'h0; // @[Mux.scala 19:72:@41623.4]
  assign _T_97568 = {_T_96971,_T_96970,_T_96969,_T_96968,_T_96967,_T_96966,_T_96965,_T_96964}; // @[Mux.scala 19:72:@41630.4]
  assign _T_97576 = {_T_96963,_T_96962,_T_96961,_T_96960,_T_96959,_T_96958,_T_96973,_T_96972,_T_97568}; // @[Mux.scala 19:72:@41638.4]
  assign _T_97578 = _T_90418 ? _T_97576 : 16'h0; // @[Mux.scala 19:72:@41639.4]
  assign _T_97585 = {_T_97042,_T_97041,_T_97040,_T_97039,_T_97038,_T_97037,_T_97036,_T_97035}; // @[Mux.scala 19:72:@41646.4]
  assign _T_97593 = {_T_97034,_T_97033,_T_97032,_T_97031,_T_97030,_T_97045,_T_97044,_T_97043,_T_97585}; // @[Mux.scala 19:72:@41654.4]
  assign _T_97595 = _T_90419 ? _T_97593 : 16'h0; // @[Mux.scala 19:72:@41655.4]
  assign _T_97602 = {_T_97113,_T_97112,_T_97111,_T_97110,_T_97109,_T_97108,_T_97107,_T_97106}; // @[Mux.scala 19:72:@41662.4]
  assign _T_97610 = {_T_97105,_T_97104,_T_97103,_T_97102,_T_97117,_T_97116,_T_97115,_T_97114,_T_97602}; // @[Mux.scala 19:72:@41670.4]
  assign _T_97612 = _T_90420 ? _T_97610 : 16'h0; // @[Mux.scala 19:72:@41671.4]
  assign _T_97619 = {_T_97184,_T_97183,_T_97182,_T_97181,_T_97180,_T_97179,_T_97178,_T_97177}; // @[Mux.scala 19:72:@41678.4]
  assign _T_97627 = {_T_97176,_T_97175,_T_97174,_T_97189,_T_97188,_T_97187,_T_97186,_T_97185,_T_97619}; // @[Mux.scala 19:72:@41686.4]
  assign _T_97629 = _T_90421 ? _T_97627 : 16'h0; // @[Mux.scala 19:72:@41687.4]
  assign _T_97636 = {_T_97255,_T_97254,_T_97253,_T_97252,_T_97251,_T_97250,_T_97249,_T_97248}; // @[Mux.scala 19:72:@41694.4]
  assign _T_97644 = {_T_97247,_T_97246,_T_97261,_T_97260,_T_97259,_T_97258,_T_97257,_T_97256,_T_97636}; // @[Mux.scala 19:72:@41702.4]
  assign _T_97646 = _T_90422 ? _T_97644 : 16'h0; // @[Mux.scala 19:72:@41703.4]
  assign _T_97653 = {_T_97326,_T_97325,_T_97324,_T_97323,_T_97322,_T_97321,_T_97320,_T_97319}; // @[Mux.scala 19:72:@41710.4]
  assign _T_97661 = {_T_97318,_T_97333,_T_97332,_T_97331,_T_97330,_T_97329,_T_97328,_T_97327,_T_97653}; // @[Mux.scala 19:72:@41718.4]
  assign _T_97663 = _T_90423 ? _T_97661 : 16'h0; // @[Mux.scala 19:72:@41719.4]
  assign _T_97664 = _T_97408 | _T_97425; // @[Mux.scala 19:72:@41720.4]
  assign _T_97665 = _T_97664 | _T_97442; // @[Mux.scala 19:72:@41721.4]
  assign _T_97666 = _T_97665 | _T_97459; // @[Mux.scala 19:72:@41722.4]
  assign _T_97667 = _T_97666 | _T_97476; // @[Mux.scala 19:72:@41723.4]
  assign _T_97668 = _T_97667 | _T_97493; // @[Mux.scala 19:72:@41724.4]
  assign _T_97669 = _T_97668 | _T_97510; // @[Mux.scala 19:72:@41725.4]
  assign _T_97670 = _T_97669 | _T_97527; // @[Mux.scala 19:72:@41726.4]
  assign _T_97671 = _T_97670 | _T_97544; // @[Mux.scala 19:72:@41727.4]
  assign _T_97672 = _T_97671 | _T_97561; // @[Mux.scala 19:72:@41728.4]
  assign _T_97673 = _T_97672 | _T_97578; // @[Mux.scala 19:72:@41729.4]
  assign _T_97674 = _T_97673 | _T_97595; // @[Mux.scala 19:72:@41730.4]
  assign _T_97675 = _T_97674 | _T_97612; // @[Mux.scala 19:72:@41731.4]
  assign _T_97676 = _T_97675 | _T_97629; // @[Mux.scala 19:72:@41732.4]
  assign _T_97677 = _T_97676 | _T_97646; // @[Mux.scala 19:72:@41733.4]
  assign _T_97678 = _T_97677 | _T_97663; // @[Mux.scala 19:72:@41734.4]
  assign outputPriorityPorts_0_0 = _T_97678[0]; // @[Mux.scala 19:72:@41738.4]
  assign outputPriorityPorts_0_1 = _T_97678[1]; // @[Mux.scala 19:72:@41740.4]
  assign outputPriorityPorts_0_2 = _T_97678[2]; // @[Mux.scala 19:72:@41742.4]
  assign outputPriorityPorts_0_3 = _T_97678[3]; // @[Mux.scala 19:72:@41744.4]
  assign outputPriorityPorts_0_4 = _T_97678[4]; // @[Mux.scala 19:72:@41746.4]
  assign outputPriorityPorts_0_5 = _T_97678[5]; // @[Mux.scala 19:72:@41748.4]
  assign outputPriorityPorts_0_6 = _T_97678[6]; // @[Mux.scala 19:72:@41750.4]
  assign outputPriorityPorts_0_7 = _T_97678[7]; // @[Mux.scala 19:72:@41752.4]
  assign outputPriorityPorts_0_8 = _T_97678[8]; // @[Mux.scala 19:72:@41754.4]
  assign outputPriorityPorts_0_9 = _T_97678[9]; // @[Mux.scala 19:72:@41756.4]
  assign outputPriorityPorts_0_10 = _T_97678[10]; // @[Mux.scala 19:72:@41758.4]
  assign outputPriorityPorts_0_11 = _T_97678[11]; // @[Mux.scala 19:72:@41760.4]
  assign outputPriorityPorts_0_12 = _T_97678[12]; // @[Mux.scala 19:72:@41762.4]
  assign outputPriorityPorts_0_13 = _T_97678[13]; // @[Mux.scala 19:72:@41764.4]
  assign outputPriorityPorts_0_14 = _T_97678[14]; // @[Mux.scala 19:72:@41766.4]
  assign outputPriorityPorts_0_15 = _T_97678[15]; // @[Mux.scala 19:72:@41768.4]
  assign _T_97822 = portQ_0 & _T_94435; // @[LoadQueue.scala 298:83:@41787.4]
  assign _T_97825 = portQ_1 & _T_94438; // @[LoadQueue.scala 298:83:@41789.4]
  assign _T_97828 = portQ_2 & _T_94441; // @[LoadQueue.scala 298:83:@41791.4]
  assign _T_97831 = portQ_3 & _T_94444; // @[LoadQueue.scala 298:83:@41793.4]
  assign _T_97834 = portQ_4 & _T_94447; // @[LoadQueue.scala 298:83:@41795.4]
  assign _T_97837 = portQ_5 & _T_94450; // @[LoadQueue.scala 298:83:@41797.4]
  assign _T_97840 = portQ_6 & _T_94453; // @[LoadQueue.scala 298:83:@41799.4]
  assign _T_97843 = portQ_7 & _T_94456; // @[LoadQueue.scala 298:83:@41801.4]
  assign _T_97846 = portQ_8 & _T_94459; // @[LoadQueue.scala 298:83:@41803.4]
  assign _T_97849 = portQ_9 & _T_94462; // @[LoadQueue.scala 298:83:@41805.4]
  assign _T_97852 = portQ_10 & _T_94465; // @[LoadQueue.scala 298:83:@41807.4]
  assign _T_97855 = portQ_11 & _T_94468; // @[LoadQueue.scala 298:83:@41809.4]
  assign _T_97858 = portQ_12 & _T_94471; // @[LoadQueue.scala 298:83:@41811.4]
  assign _T_97861 = portQ_13 & _T_94474; // @[LoadQueue.scala 298:83:@41813.4]
  assign _T_97864 = portQ_14 & _T_94477; // @[LoadQueue.scala 298:83:@41815.4]
  assign _T_97867 = portQ_15 & _T_94480; // @[LoadQueue.scala 298:83:@41817.4]
  assign _T_97950 = _T_97867 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41871.4]
  assign _T_97951 = _T_97864 ? 16'h4000 : _T_97950; // @[Mux.scala 31:69:@41872.4]
  assign _T_97952 = _T_97861 ? 16'h2000 : _T_97951; // @[Mux.scala 31:69:@41873.4]
  assign _T_97953 = _T_97858 ? 16'h1000 : _T_97952; // @[Mux.scala 31:69:@41874.4]
  assign _T_97954 = _T_97855 ? 16'h800 : _T_97953; // @[Mux.scala 31:69:@41875.4]
  assign _T_97955 = _T_97852 ? 16'h400 : _T_97954; // @[Mux.scala 31:69:@41876.4]
  assign _T_97956 = _T_97849 ? 16'h200 : _T_97955; // @[Mux.scala 31:69:@41877.4]
  assign _T_97957 = _T_97846 ? 16'h100 : _T_97956; // @[Mux.scala 31:69:@41878.4]
  assign _T_97958 = _T_97843 ? 16'h80 : _T_97957; // @[Mux.scala 31:69:@41879.4]
  assign _T_97959 = _T_97840 ? 16'h40 : _T_97958; // @[Mux.scala 31:69:@41880.4]
  assign _T_97960 = _T_97837 ? 16'h20 : _T_97959; // @[Mux.scala 31:69:@41881.4]
  assign _T_97961 = _T_97834 ? 16'h10 : _T_97960; // @[Mux.scala 31:69:@41882.4]
  assign _T_97962 = _T_97831 ? 16'h8 : _T_97961; // @[Mux.scala 31:69:@41883.4]
  assign _T_97963 = _T_97828 ? 16'h4 : _T_97962; // @[Mux.scala 31:69:@41884.4]
  assign _T_97964 = _T_97825 ? 16'h2 : _T_97963; // @[Mux.scala 31:69:@41885.4]
  assign _T_97965 = _T_97822 ? 16'h1 : _T_97964; // @[Mux.scala 31:69:@41886.4]
  assign _T_97966 = _T_97965[0]; // @[OneHot.scala 66:30:@41887.4]
  assign _T_97967 = _T_97965[1]; // @[OneHot.scala 66:30:@41888.4]
  assign _T_97968 = _T_97965[2]; // @[OneHot.scala 66:30:@41889.4]
  assign _T_97969 = _T_97965[3]; // @[OneHot.scala 66:30:@41890.4]
  assign _T_97970 = _T_97965[4]; // @[OneHot.scala 66:30:@41891.4]
  assign _T_97971 = _T_97965[5]; // @[OneHot.scala 66:30:@41892.4]
  assign _T_97972 = _T_97965[6]; // @[OneHot.scala 66:30:@41893.4]
  assign _T_97973 = _T_97965[7]; // @[OneHot.scala 66:30:@41894.4]
  assign _T_97974 = _T_97965[8]; // @[OneHot.scala 66:30:@41895.4]
  assign _T_97975 = _T_97965[9]; // @[OneHot.scala 66:30:@41896.4]
  assign _T_97976 = _T_97965[10]; // @[OneHot.scala 66:30:@41897.4]
  assign _T_97977 = _T_97965[11]; // @[OneHot.scala 66:30:@41898.4]
  assign _T_97978 = _T_97965[12]; // @[OneHot.scala 66:30:@41899.4]
  assign _T_97979 = _T_97965[13]; // @[OneHot.scala 66:30:@41900.4]
  assign _T_97980 = _T_97965[14]; // @[OneHot.scala 66:30:@41901.4]
  assign _T_97981 = _T_97965[15]; // @[OneHot.scala 66:30:@41902.4]
  assign _T_98022 = _T_97822 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41920.4]
  assign _T_98023 = _T_97867 ? 16'h4000 : _T_98022; // @[Mux.scala 31:69:@41921.4]
  assign _T_98024 = _T_97864 ? 16'h2000 : _T_98023; // @[Mux.scala 31:69:@41922.4]
  assign _T_98025 = _T_97861 ? 16'h1000 : _T_98024; // @[Mux.scala 31:69:@41923.4]
  assign _T_98026 = _T_97858 ? 16'h800 : _T_98025; // @[Mux.scala 31:69:@41924.4]
  assign _T_98027 = _T_97855 ? 16'h400 : _T_98026; // @[Mux.scala 31:69:@41925.4]
  assign _T_98028 = _T_97852 ? 16'h200 : _T_98027; // @[Mux.scala 31:69:@41926.4]
  assign _T_98029 = _T_97849 ? 16'h100 : _T_98028; // @[Mux.scala 31:69:@41927.4]
  assign _T_98030 = _T_97846 ? 16'h80 : _T_98029; // @[Mux.scala 31:69:@41928.4]
  assign _T_98031 = _T_97843 ? 16'h40 : _T_98030; // @[Mux.scala 31:69:@41929.4]
  assign _T_98032 = _T_97840 ? 16'h20 : _T_98031; // @[Mux.scala 31:69:@41930.4]
  assign _T_98033 = _T_97837 ? 16'h10 : _T_98032; // @[Mux.scala 31:69:@41931.4]
  assign _T_98034 = _T_97834 ? 16'h8 : _T_98033; // @[Mux.scala 31:69:@41932.4]
  assign _T_98035 = _T_97831 ? 16'h4 : _T_98034; // @[Mux.scala 31:69:@41933.4]
  assign _T_98036 = _T_97828 ? 16'h2 : _T_98035; // @[Mux.scala 31:69:@41934.4]
  assign _T_98037 = _T_97825 ? 16'h1 : _T_98036; // @[Mux.scala 31:69:@41935.4]
  assign _T_98038 = _T_98037[0]; // @[OneHot.scala 66:30:@41936.4]
  assign _T_98039 = _T_98037[1]; // @[OneHot.scala 66:30:@41937.4]
  assign _T_98040 = _T_98037[2]; // @[OneHot.scala 66:30:@41938.4]
  assign _T_98041 = _T_98037[3]; // @[OneHot.scala 66:30:@41939.4]
  assign _T_98042 = _T_98037[4]; // @[OneHot.scala 66:30:@41940.4]
  assign _T_98043 = _T_98037[5]; // @[OneHot.scala 66:30:@41941.4]
  assign _T_98044 = _T_98037[6]; // @[OneHot.scala 66:30:@41942.4]
  assign _T_98045 = _T_98037[7]; // @[OneHot.scala 66:30:@41943.4]
  assign _T_98046 = _T_98037[8]; // @[OneHot.scala 66:30:@41944.4]
  assign _T_98047 = _T_98037[9]; // @[OneHot.scala 66:30:@41945.4]
  assign _T_98048 = _T_98037[10]; // @[OneHot.scala 66:30:@41946.4]
  assign _T_98049 = _T_98037[11]; // @[OneHot.scala 66:30:@41947.4]
  assign _T_98050 = _T_98037[12]; // @[OneHot.scala 66:30:@41948.4]
  assign _T_98051 = _T_98037[13]; // @[OneHot.scala 66:30:@41949.4]
  assign _T_98052 = _T_98037[14]; // @[OneHot.scala 66:30:@41950.4]
  assign _T_98053 = _T_98037[15]; // @[OneHot.scala 66:30:@41951.4]
  assign _T_98094 = _T_97825 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41969.4]
  assign _T_98095 = _T_97822 ? 16'h4000 : _T_98094; // @[Mux.scala 31:69:@41970.4]
  assign _T_98096 = _T_97867 ? 16'h2000 : _T_98095; // @[Mux.scala 31:69:@41971.4]
  assign _T_98097 = _T_97864 ? 16'h1000 : _T_98096; // @[Mux.scala 31:69:@41972.4]
  assign _T_98098 = _T_97861 ? 16'h800 : _T_98097; // @[Mux.scala 31:69:@41973.4]
  assign _T_98099 = _T_97858 ? 16'h400 : _T_98098; // @[Mux.scala 31:69:@41974.4]
  assign _T_98100 = _T_97855 ? 16'h200 : _T_98099; // @[Mux.scala 31:69:@41975.4]
  assign _T_98101 = _T_97852 ? 16'h100 : _T_98100; // @[Mux.scala 31:69:@41976.4]
  assign _T_98102 = _T_97849 ? 16'h80 : _T_98101; // @[Mux.scala 31:69:@41977.4]
  assign _T_98103 = _T_97846 ? 16'h40 : _T_98102; // @[Mux.scala 31:69:@41978.4]
  assign _T_98104 = _T_97843 ? 16'h20 : _T_98103; // @[Mux.scala 31:69:@41979.4]
  assign _T_98105 = _T_97840 ? 16'h10 : _T_98104; // @[Mux.scala 31:69:@41980.4]
  assign _T_98106 = _T_97837 ? 16'h8 : _T_98105; // @[Mux.scala 31:69:@41981.4]
  assign _T_98107 = _T_97834 ? 16'h4 : _T_98106; // @[Mux.scala 31:69:@41982.4]
  assign _T_98108 = _T_97831 ? 16'h2 : _T_98107; // @[Mux.scala 31:69:@41983.4]
  assign _T_98109 = _T_97828 ? 16'h1 : _T_98108; // @[Mux.scala 31:69:@41984.4]
  assign _T_98110 = _T_98109[0]; // @[OneHot.scala 66:30:@41985.4]
  assign _T_98111 = _T_98109[1]; // @[OneHot.scala 66:30:@41986.4]
  assign _T_98112 = _T_98109[2]; // @[OneHot.scala 66:30:@41987.4]
  assign _T_98113 = _T_98109[3]; // @[OneHot.scala 66:30:@41988.4]
  assign _T_98114 = _T_98109[4]; // @[OneHot.scala 66:30:@41989.4]
  assign _T_98115 = _T_98109[5]; // @[OneHot.scala 66:30:@41990.4]
  assign _T_98116 = _T_98109[6]; // @[OneHot.scala 66:30:@41991.4]
  assign _T_98117 = _T_98109[7]; // @[OneHot.scala 66:30:@41992.4]
  assign _T_98118 = _T_98109[8]; // @[OneHot.scala 66:30:@41993.4]
  assign _T_98119 = _T_98109[9]; // @[OneHot.scala 66:30:@41994.4]
  assign _T_98120 = _T_98109[10]; // @[OneHot.scala 66:30:@41995.4]
  assign _T_98121 = _T_98109[11]; // @[OneHot.scala 66:30:@41996.4]
  assign _T_98122 = _T_98109[12]; // @[OneHot.scala 66:30:@41997.4]
  assign _T_98123 = _T_98109[13]; // @[OneHot.scala 66:30:@41998.4]
  assign _T_98124 = _T_98109[14]; // @[OneHot.scala 66:30:@41999.4]
  assign _T_98125 = _T_98109[15]; // @[OneHot.scala 66:30:@42000.4]
  assign _T_98166 = _T_97828 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42018.4]
  assign _T_98167 = _T_97825 ? 16'h4000 : _T_98166; // @[Mux.scala 31:69:@42019.4]
  assign _T_98168 = _T_97822 ? 16'h2000 : _T_98167; // @[Mux.scala 31:69:@42020.4]
  assign _T_98169 = _T_97867 ? 16'h1000 : _T_98168; // @[Mux.scala 31:69:@42021.4]
  assign _T_98170 = _T_97864 ? 16'h800 : _T_98169; // @[Mux.scala 31:69:@42022.4]
  assign _T_98171 = _T_97861 ? 16'h400 : _T_98170; // @[Mux.scala 31:69:@42023.4]
  assign _T_98172 = _T_97858 ? 16'h200 : _T_98171; // @[Mux.scala 31:69:@42024.4]
  assign _T_98173 = _T_97855 ? 16'h100 : _T_98172; // @[Mux.scala 31:69:@42025.4]
  assign _T_98174 = _T_97852 ? 16'h80 : _T_98173; // @[Mux.scala 31:69:@42026.4]
  assign _T_98175 = _T_97849 ? 16'h40 : _T_98174; // @[Mux.scala 31:69:@42027.4]
  assign _T_98176 = _T_97846 ? 16'h20 : _T_98175; // @[Mux.scala 31:69:@42028.4]
  assign _T_98177 = _T_97843 ? 16'h10 : _T_98176; // @[Mux.scala 31:69:@42029.4]
  assign _T_98178 = _T_97840 ? 16'h8 : _T_98177; // @[Mux.scala 31:69:@42030.4]
  assign _T_98179 = _T_97837 ? 16'h4 : _T_98178; // @[Mux.scala 31:69:@42031.4]
  assign _T_98180 = _T_97834 ? 16'h2 : _T_98179; // @[Mux.scala 31:69:@42032.4]
  assign _T_98181 = _T_97831 ? 16'h1 : _T_98180; // @[Mux.scala 31:69:@42033.4]
  assign _T_98182 = _T_98181[0]; // @[OneHot.scala 66:30:@42034.4]
  assign _T_98183 = _T_98181[1]; // @[OneHot.scala 66:30:@42035.4]
  assign _T_98184 = _T_98181[2]; // @[OneHot.scala 66:30:@42036.4]
  assign _T_98185 = _T_98181[3]; // @[OneHot.scala 66:30:@42037.4]
  assign _T_98186 = _T_98181[4]; // @[OneHot.scala 66:30:@42038.4]
  assign _T_98187 = _T_98181[5]; // @[OneHot.scala 66:30:@42039.4]
  assign _T_98188 = _T_98181[6]; // @[OneHot.scala 66:30:@42040.4]
  assign _T_98189 = _T_98181[7]; // @[OneHot.scala 66:30:@42041.4]
  assign _T_98190 = _T_98181[8]; // @[OneHot.scala 66:30:@42042.4]
  assign _T_98191 = _T_98181[9]; // @[OneHot.scala 66:30:@42043.4]
  assign _T_98192 = _T_98181[10]; // @[OneHot.scala 66:30:@42044.4]
  assign _T_98193 = _T_98181[11]; // @[OneHot.scala 66:30:@42045.4]
  assign _T_98194 = _T_98181[12]; // @[OneHot.scala 66:30:@42046.4]
  assign _T_98195 = _T_98181[13]; // @[OneHot.scala 66:30:@42047.4]
  assign _T_98196 = _T_98181[14]; // @[OneHot.scala 66:30:@42048.4]
  assign _T_98197 = _T_98181[15]; // @[OneHot.scala 66:30:@42049.4]
  assign _T_98238 = _T_97831 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42067.4]
  assign _T_98239 = _T_97828 ? 16'h4000 : _T_98238; // @[Mux.scala 31:69:@42068.4]
  assign _T_98240 = _T_97825 ? 16'h2000 : _T_98239; // @[Mux.scala 31:69:@42069.4]
  assign _T_98241 = _T_97822 ? 16'h1000 : _T_98240; // @[Mux.scala 31:69:@42070.4]
  assign _T_98242 = _T_97867 ? 16'h800 : _T_98241; // @[Mux.scala 31:69:@42071.4]
  assign _T_98243 = _T_97864 ? 16'h400 : _T_98242; // @[Mux.scala 31:69:@42072.4]
  assign _T_98244 = _T_97861 ? 16'h200 : _T_98243; // @[Mux.scala 31:69:@42073.4]
  assign _T_98245 = _T_97858 ? 16'h100 : _T_98244; // @[Mux.scala 31:69:@42074.4]
  assign _T_98246 = _T_97855 ? 16'h80 : _T_98245; // @[Mux.scala 31:69:@42075.4]
  assign _T_98247 = _T_97852 ? 16'h40 : _T_98246; // @[Mux.scala 31:69:@42076.4]
  assign _T_98248 = _T_97849 ? 16'h20 : _T_98247; // @[Mux.scala 31:69:@42077.4]
  assign _T_98249 = _T_97846 ? 16'h10 : _T_98248; // @[Mux.scala 31:69:@42078.4]
  assign _T_98250 = _T_97843 ? 16'h8 : _T_98249; // @[Mux.scala 31:69:@42079.4]
  assign _T_98251 = _T_97840 ? 16'h4 : _T_98250; // @[Mux.scala 31:69:@42080.4]
  assign _T_98252 = _T_97837 ? 16'h2 : _T_98251; // @[Mux.scala 31:69:@42081.4]
  assign _T_98253 = _T_97834 ? 16'h1 : _T_98252; // @[Mux.scala 31:69:@42082.4]
  assign _T_98254 = _T_98253[0]; // @[OneHot.scala 66:30:@42083.4]
  assign _T_98255 = _T_98253[1]; // @[OneHot.scala 66:30:@42084.4]
  assign _T_98256 = _T_98253[2]; // @[OneHot.scala 66:30:@42085.4]
  assign _T_98257 = _T_98253[3]; // @[OneHot.scala 66:30:@42086.4]
  assign _T_98258 = _T_98253[4]; // @[OneHot.scala 66:30:@42087.4]
  assign _T_98259 = _T_98253[5]; // @[OneHot.scala 66:30:@42088.4]
  assign _T_98260 = _T_98253[6]; // @[OneHot.scala 66:30:@42089.4]
  assign _T_98261 = _T_98253[7]; // @[OneHot.scala 66:30:@42090.4]
  assign _T_98262 = _T_98253[8]; // @[OneHot.scala 66:30:@42091.4]
  assign _T_98263 = _T_98253[9]; // @[OneHot.scala 66:30:@42092.4]
  assign _T_98264 = _T_98253[10]; // @[OneHot.scala 66:30:@42093.4]
  assign _T_98265 = _T_98253[11]; // @[OneHot.scala 66:30:@42094.4]
  assign _T_98266 = _T_98253[12]; // @[OneHot.scala 66:30:@42095.4]
  assign _T_98267 = _T_98253[13]; // @[OneHot.scala 66:30:@42096.4]
  assign _T_98268 = _T_98253[14]; // @[OneHot.scala 66:30:@42097.4]
  assign _T_98269 = _T_98253[15]; // @[OneHot.scala 66:30:@42098.4]
  assign _T_98310 = _T_97834 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42116.4]
  assign _T_98311 = _T_97831 ? 16'h4000 : _T_98310; // @[Mux.scala 31:69:@42117.4]
  assign _T_98312 = _T_97828 ? 16'h2000 : _T_98311; // @[Mux.scala 31:69:@42118.4]
  assign _T_98313 = _T_97825 ? 16'h1000 : _T_98312; // @[Mux.scala 31:69:@42119.4]
  assign _T_98314 = _T_97822 ? 16'h800 : _T_98313; // @[Mux.scala 31:69:@42120.4]
  assign _T_98315 = _T_97867 ? 16'h400 : _T_98314; // @[Mux.scala 31:69:@42121.4]
  assign _T_98316 = _T_97864 ? 16'h200 : _T_98315; // @[Mux.scala 31:69:@42122.4]
  assign _T_98317 = _T_97861 ? 16'h100 : _T_98316; // @[Mux.scala 31:69:@42123.4]
  assign _T_98318 = _T_97858 ? 16'h80 : _T_98317; // @[Mux.scala 31:69:@42124.4]
  assign _T_98319 = _T_97855 ? 16'h40 : _T_98318; // @[Mux.scala 31:69:@42125.4]
  assign _T_98320 = _T_97852 ? 16'h20 : _T_98319; // @[Mux.scala 31:69:@42126.4]
  assign _T_98321 = _T_97849 ? 16'h10 : _T_98320; // @[Mux.scala 31:69:@42127.4]
  assign _T_98322 = _T_97846 ? 16'h8 : _T_98321; // @[Mux.scala 31:69:@42128.4]
  assign _T_98323 = _T_97843 ? 16'h4 : _T_98322; // @[Mux.scala 31:69:@42129.4]
  assign _T_98324 = _T_97840 ? 16'h2 : _T_98323; // @[Mux.scala 31:69:@42130.4]
  assign _T_98325 = _T_97837 ? 16'h1 : _T_98324; // @[Mux.scala 31:69:@42131.4]
  assign _T_98326 = _T_98325[0]; // @[OneHot.scala 66:30:@42132.4]
  assign _T_98327 = _T_98325[1]; // @[OneHot.scala 66:30:@42133.4]
  assign _T_98328 = _T_98325[2]; // @[OneHot.scala 66:30:@42134.4]
  assign _T_98329 = _T_98325[3]; // @[OneHot.scala 66:30:@42135.4]
  assign _T_98330 = _T_98325[4]; // @[OneHot.scala 66:30:@42136.4]
  assign _T_98331 = _T_98325[5]; // @[OneHot.scala 66:30:@42137.4]
  assign _T_98332 = _T_98325[6]; // @[OneHot.scala 66:30:@42138.4]
  assign _T_98333 = _T_98325[7]; // @[OneHot.scala 66:30:@42139.4]
  assign _T_98334 = _T_98325[8]; // @[OneHot.scala 66:30:@42140.4]
  assign _T_98335 = _T_98325[9]; // @[OneHot.scala 66:30:@42141.4]
  assign _T_98336 = _T_98325[10]; // @[OneHot.scala 66:30:@42142.4]
  assign _T_98337 = _T_98325[11]; // @[OneHot.scala 66:30:@42143.4]
  assign _T_98338 = _T_98325[12]; // @[OneHot.scala 66:30:@42144.4]
  assign _T_98339 = _T_98325[13]; // @[OneHot.scala 66:30:@42145.4]
  assign _T_98340 = _T_98325[14]; // @[OneHot.scala 66:30:@42146.4]
  assign _T_98341 = _T_98325[15]; // @[OneHot.scala 66:30:@42147.4]
  assign _T_98382 = _T_97837 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42165.4]
  assign _T_98383 = _T_97834 ? 16'h4000 : _T_98382; // @[Mux.scala 31:69:@42166.4]
  assign _T_98384 = _T_97831 ? 16'h2000 : _T_98383; // @[Mux.scala 31:69:@42167.4]
  assign _T_98385 = _T_97828 ? 16'h1000 : _T_98384; // @[Mux.scala 31:69:@42168.4]
  assign _T_98386 = _T_97825 ? 16'h800 : _T_98385; // @[Mux.scala 31:69:@42169.4]
  assign _T_98387 = _T_97822 ? 16'h400 : _T_98386; // @[Mux.scala 31:69:@42170.4]
  assign _T_98388 = _T_97867 ? 16'h200 : _T_98387; // @[Mux.scala 31:69:@42171.4]
  assign _T_98389 = _T_97864 ? 16'h100 : _T_98388; // @[Mux.scala 31:69:@42172.4]
  assign _T_98390 = _T_97861 ? 16'h80 : _T_98389; // @[Mux.scala 31:69:@42173.4]
  assign _T_98391 = _T_97858 ? 16'h40 : _T_98390; // @[Mux.scala 31:69:@42174.4]
  assign _T_98392 = _T_97855 ? 16'h20 : _T_98391; // @[Mux.scala 31:69:@42175.4]
  assign _T_98393 = _T_97852 ? 16'h10 : _T_98392; // @[Mux.scala 31:69:@42176.4]
  assign _T_98394 = _T_97849 ? 16'h8 : _T_98393; // @[Mux.scala 31:69:@42177.4]
  assign _T_98395 = _T_97846 ? 16'h4 : _T_98394; // @[Mux.scala 31:69:@42178.4]
  assign _T_98396 = _T_97843 ? 16'h2 : _T_98395; // @[Mux.scala 31:69:@42179.4]
  assign _T_98397 = _T_97840 ? 16'h1 : _T_98396; // @[Mux.scala 31:69:@42180.4]
  assign _T_98398 = _T_98397[0]; // @[OneHot.scala 66:30:@42181.4]
  assign _T_98399 = _T_98397[1]; // @[OneHot.scala 66:30:@42182.4]
  assign _T_98400 = _T_98397[2]; // @[OneHot.scala 66:30:@42183.4]
  assign _T_98401 = _T_98397[3]; // @[OneHot.scala 66:30:@42184.4]
  assign _T_98402 = _T_98397[4]; // @[OneHot.scala 66:30:@42185.4]
  assign _T_98403 = _T_98397[5]; // @[OneHot.scala 66:30:@42186.4]
  assign _T_98404 = _T_98397[6]; // @[OneHot.scala 66:30:@42187.4]
  assign _T_98405 = _T_98397[7]; // @[OneHot.scala 66:30:@42188.4]
  assign _T_98406 = _T_98397[8]; // @[OneHot.scala 66:30:@42189.4]
  assign _T_98407 = _T_98397[9]; // @[OneHot.scala 66:30:@42190.4]
  assign _T_98408 = _T_98397[10]; // @[OneHot.scala 66:30:@42191.4]
  assign _T_98409 = _T_98397[11]; // @[OneHot.scala 66:30:@42192.4]
  assign _T_98410 = _T_98397[12]; // @[OneHot.scala 66:30:@42193.4]
  assign _T_98411 = _T_98397[13]; // @[OneHot.scala 66:30:@42194.4]
  assign _T_98412 = _T_98397[14]; // @[OneHot.scala 66:30:@42195.4]
  assign _T_98413 = _T_98397[15]; // @[OneHot.scala 66:30:@42196.4]
  assign _T_98454 = _T_97840 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42214.4]
  assign _T_98455 = _T_97837 ? 16'h4000 : _T_98454; // @[Mux.scala 31:69:@42215.4]
  assign _T_98456 = _T_97834 ? 16'h2000 : _T_98455; // @[Mux.scala 31:69:@42216.4]
  assign _T_98457 = _T_97831 ? 16'h1000 : _T_98456; // @[Mux.scala 31:69:@42217.4]
  assign _T_98458 = _T_97828 ? 16'h800 : _T_98457; // @[Mux.scala 31:69:@42218.4]
  assign _T_98459 = _T_97825 ? 16'h400 : _T_98458; // @[Mux.scala 31:69:@42219.4]
  assign _T_98460 = _T_97822 ? 16'h200 : _T_98459; // @[Mux.scala 31:69:@42220.4]
  assign _T_98461 = _T_97867 ? 16'h100 : _T_98460; // @[Mux.scala 31:69:@42221.4]
  assign _T_98462 = _T_97864 ? 16'h80 : _T_98461; // @[Mux.scala 31:69:@42222.4]
  assign _T_98463 = _T_97861 ? 16'h40 : _T_98462; // @[Mux.scala 31:69:@42223.4]
  assign _T_98464 = _T_97858 ? 16'h20 : _T_98463; // @[Mux.scala 31:69:@42224.4]
  assign _T_98465 = _T_97855 ? 16'h10 : _T_98464; // @[Mux.scala 31:69:@42225.4]
  assign _T_98466 = _T_97852 ? 16'h8 : _T_98465; // @[Mux.scala 31:69:@42226.4]
  assign _T_98467 = _T_97849 ? 16'h4 : _T_98466; // @[Mux.scala 31:69:@42227.4]
  assign _T_98468 = _T_97846 ? 16'h2 : _T_98467; // @[Mux.scala 31:69:@42228.4]
  assign _T_98469 = _T_97843 ? 16'h1 : _T_98468; // @[Mux.scala 31:69:@42229.4]
  assign _T_98470 = _T_98469[0]; // @[OneHot.scala 66:30:@42230.4]
  assign _T_98471 = _T_98469[1]; // @[OneHot.scala 66:30:@42231.4]
  assign _T_98472 = _T_98469[2]; // @[OneHot.scala 66:30:@42232.4]
  assign _T_98473 = _T_98469[3]; // @[OneHot.scala 66:30:@42233.4]
  assign _T_98474 = _T_98469[4]; // @[OneHot.scala 66:30:@42234.4]
  assign _T_98475 = _T_98469[5]; // @[OneHot.scala 66:30:@42235.4]
  assign _T_98476 = _T_98469[6]; // @[OneHot.scala 66:30:@42236.4]
  assign _T_98477 = _T_98469[7]; // @[OneHot.scala 66:30:@42237.4]
  assign _T_98478 = _T_98469[8]; // @[OneHot.scala 66:30:@42238.4]
  assign _T_98479 = _T_98469[9]; // @[OneHot.scala 66:30:@42239.4]
  assign _T_98480 = _T_98469[10]; // @[OneHot.scala 66:30:@42240.4]
  assign _T_98481 = _T_98469[11]; // @[OneHot.scala 66:30:@42241.4]
  assign _T_98482 = _T_98469[12]; // @[OneHot.scala 66:30:@42242.4]
  assign _T_98483 = _T_98469[13]; // @[OneHot.scala 66:30:@42243.4]
  assign _T_98484 = _T_98469[14]; // @[OneHot.scala 66:30:@42244.4]
  assign _T_98485 = _T_98469[15]; // @[OneHot.scala 66:30:@42245.4]
  assign _T_98526 = _T_97843 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42263.4]
  assign _T_98527 = _T_97840 ? 16'h4000 : _T_98526; // @[Mux.scala 31:69:@42264.4]
  assign _T_98528 = _T_97837 ? 16'h2000 : _T_98527; // @[Mux.scala 31:69:@42265.4]
  assign _T_98529 = _T_97834 ? 16'h1000 : _T_98528; // @[Mux.scala 31:69:@42266.4]
  assign _T_98530 = _T_97831 ? 16'h800 : _T_98529; // @[Mux.scala 31:69:@42267.4]
  assign _T_98531 = _T_97828 ? 16'h400 : _T_98530; // @[Mux.scala 31:69:@42268.4]
  assign _T_98532 = _T_97825 ? 16'h200 : _T_98531; // @[Mux.scala 31:69:@42269.4]
  assign _T_98533 = _T_97822 ? 16'h100 : _T_98532; // @[Mux.scala 31:69:@42270.4]
  assign _T_98534 = _T_97867 ? 16'h80 : _T_98533; // @[Mux.scala 31:69:@42271.4]
  assign _T_98535 = _T_97864 ? 16'h40 : _T_98534; // @[Mux.scala 31:69:@42272.4]
  assign _T_98536 = _T_97861 ? 16'h20 : _T_98535; // @[Mux.scala 31:69:@42273.4]
  assign _T_98537 = _T_97858 ? 16'h10 : _T_98536; // @[Mux.scala 31:69:@42274.4]
  assign _T_98538 = _T_97855 ? 16'h8 : _T_98537; // @[Mux.scala 31:69:@42275.4]
  assign _T_98539 = _T_97852 ? 16'h4 : _T_98538; // @[Mux.scala 31:69:@42276.4]
  assign _T_98540 = _T_97849 ? 16'h2 : _T_98539; // @[Mux.scala 31:69:@42277.4]
  assign _T_98541 = _T_97846 ? 16'h1 : _T_98540; // @[Mux.scala 31:69:@42278.4]
  assign _T_98542 = _T_98541[0]; // @[OneHot.scala 66:30:@42279.4]
  assign _T_98543 = _T_98541[1]; // @[OneHot.scala 66:30:@42280.4]
  assign _T_98544 = _T_98541[2]; // @[OneHot.scala 66:30:@42281.4]
  assign _T_98545 = _T_98541[3]; // @[OneHot.scala 66:30:@42282.4]
  assign _T_98546 = _T_98541[4]; // @[OneHot.scala 66:30:@42283.4]
  assign _T_98547 = _T_98541[5]; // @[OneHot.scala 66:30:@42284.4]
  assign _T_98548 = _T_98541[6]; // @[OneHot.scala 66:30:@42285.4]
  assign _T_98549 = _T_98541[7]; // @[OneHot.scala 66:30:@42286.4]
  assign _T_98550 = _T_98541[8]; // @[OneHot.scala 66:30:@42287.4]
  assign _T_98551 = _T_98541[9]; // @[OneHot.scala 66:30:@42288.4]
  assign _T_98552 = _T_98541[10]; // @[OneHot.scala 66:30:@42289.4]
  assign _T_98553 = _T_98541[11]; // @[OneHot.scala 66:30:@42290.4]
  assign _T_98554 = _T_98541[12]; // @[OneHot.scala 66:30:@42291.4]
  assign _T_98555 = _T_98541[13]; // @[OneHot.scala 66:30:@42292.4]
  assign _T_98556 = _T_98541[14]; // @[OneHot.scala 66:30:@42293.4]
  assign _T_98557 = _T_98541[15]; // @[OneHot.scala 66:30:@42294.4]
  assign _T_98598 = _T_97846 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42312.4]
  assign _T_98599 = _T_97843 ? 16'h4000 : _T_98598; // @[Mux.scala 31:69:@42313.4]
  assign _T_98600 = _T_97840 ? 16'h2000 : _T_98599; // @[Mux.scala 31:69:@42314.4]
  assign _T_98601 = _T_97837 ? 16'h1000 : _T_98600; // @[Mux.scala 31:69:@42315.4]
  assign _T_98602 = _T_97834 ? 16'h800 : _T_98601; // @[Mux.scala 31:69:@42316.4]
  assign _T_98603 = _T_97831 ? 16'h400 : _T_98602; // @[Mux.scala 31:69:@42317.4]
  assign _T_98604 = _T_97828 ? 16'h200 : _T_98603; // @[Mux.scala 31:69:@42318.4]
  assign _T_98605 = _T_97825 ? 16'h100 : _T_98604; // @[Mux.scala 31:69:@42319.4]
  assign _T_98606 = _T_97822 ? 16'h80 : _T_98605; // @[Mux.scala 31:69:@42320.4]
  assign _T_98607 = _T_97867 ? 16'h40 : _T_98606; // @[Mux.scala 31:69:@42321.4]
  assign _T_98608 = _T_97864 ? 16'h20 : _T_98607; // @[Mux.scala 31:69:@42322.4]
  assign _T_98609 = _T_97861 ? 16'h10 : _T_98608; // @[Mux.scala 31:69:@42323.4]
  assign _T_98610 = _T_97858 ? 16'h8 : _T_98609; // @[Mux.scala 31:69:@42324.4]
  assign _T_98611 = _T_97855 ? 16'h4 : _T_98610; // @[Mux.scala 31:69:@42325.4]
  assign _T_98612 = _T_97852 ? 16'h2 : _T_98611; // @[Mux.scala 31:69:@42326.4]
  assign _T_98613 = _T_97849 ? 16'h1 : _T_98612; // @[Mux.scala 31:69:@42327.4]
  assign _T_98614 = _T_98613[0]; // @[OneHot.scala 66:30:@42328.4]
  assign _T_98615 = _T_98613[1]; // @[OneHot.scala 66:30:@42329.4]
  assign _T_98616 = _T_98613[2]; // @[OneHot.scala 66:30:@42330.4]
  assign _T_98617 = _T_98613[3]; // @[OneHot.scala 66:30:@42331.4]
  assign _T_98618 = _T_98613[4]; // @[OneHot.scala 66:30:@42332.4]
  assign _T_98619 = _T_98613[5]; // @[OneHot.scala 66:30:@42333.4]
  assign _T_98620 = _T_98613[6]; // @[OneHot.scala 66:30:@42334.4]
  assign _T_98621 = _T_98613[7]; // @[OneHot.scala 66:30:@42335.4]
  assign _T_98622 = _T_98613[8]; // @[OneHot.scala 66:30:@42336.4]
  assign _T_98623 = _T_98613[9]; // @[OneHot.scala 66:30:@42337.4]
  assign _T_98624 = _T_98613[10]; // @[OneHot.scala 66:30:@42338.4]
  assign _T_98625 = _T_98613[11]; // @[OneHot.scala 66:30:@42339.4]
  assign _T_98626 = _T_98613[12]; // @[OneHot.scala 66:30:@42340.4]
  assign _T_98627 = _T_98613[13]; // @[OneHot.scala 66:30:@42341.4]
  assign _T_98628 = _T_98613[14]; // @[OneHot.scala 66:30:@42342.4]
  assign _T_98629 = _T_98613[15]; // @[OneHot.scala 66:30:@42343.4]
  assign _T_98670 = _T_97849 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42361.4]
  assign _T_98671 = _T_97846 ? 16'h4000 : _T_98670; // @[Mux.scala 31:69:@42362.4]
  assign _T_98672 = _T_97843 ? 16'h2000 : _T_98671; // @[Mux.scala 31:69:@42363.4]
  assign _T_98673 = _T_97840 ? 16'h1000 : _T_98672; // @[Mux.scala 31:69:@42364.4]
  assign _T_98674 = _T_97837 ? 16'h800 : _T_98673; // @[Mux.scala 31:69:@42365.4]
  assign _T_98675 = _T_97834 ? 16'h400 : _T_98674; // @[Mux.scala 31:69:@42366.4]
  assign _T_98676 = _T_97831 ? 16'h200 : _T_98675; // @[Mux.scala 31:69:@42367.4]
  assign _T_98677 = _T_97828 ? 16'h100 : _T_98676; // @[Mux.scala 31:69:@42368.4]
  assign _T_98678 = _T_97825 ? 16'h80 : _T_98677; // @[Mux.scala 31:69:@42369.4]
  assign _T_98679 = _T_97822 ? 16'h40 : _T_98678; // @[Mux.scala 31:69:@42370.4]
  assign _T_98680 = _T_97867 ? 16'h20 : _T_98679; // @[Mux.scala 31:69:@42371.4]
  assign _T_98681 = _T_97864 ? 16'h10 : _T_98680; // @[Mux.scala 31:69:@42372.4]
  assign _T_98682 = _T_97861 ? 16'h8 : _T_98681; // @[Mux.scala 31:69:@42373.4]
  assign _T_98683 = _T_97858 ? 16'h4 : _T_98682; // @[Mux.scala 31:69:@42374.4]
  assign _T_98684 = _T_97855 ? 16'h2 : _T_98683; // @[Mux.scala 31:69:@42375.4]
  assign _T_98685 = _T_97852 ? 16'h1 : _T_98684; // @[Mux.scala 31:69:@42376.4]
  assign _T_98686 = _T_98685[0]; // @[OneHot.scala 66:30:@42377.4]
  assign _T_98687 = _T_98685[1]; // @[OneHot.scala 66:30:@42378.4]
  assign _T_98688 = _T_98685[2]; // @[OneHot.scala 66:30:@42379.4]
  assign _T_98689 = _T_98685[3]; // @[OneHot.scala 66:30:@42380.4]
  assign _T_98690 = _T_98685[4]; // @[OneHot.scala 66:30:@42381.4]
  assign _T_98691 = _T_98685[5]; // @[OneHot.scala 66:30:@42382.4]
  assign _T_98692 = _T_98685[6]; // @[OneHot.scala 66:30:@42383.4]
  assign _T_98693 = _T_98685[7]; // @[OneHot.scala 66:30:@42384.4]
  assign _T_98694 = _T_98685[8]; // @[OneHot.scala 66:30:@42385.4]
  assign _T_98695 = _T_98685[9]; // @[OneHot.scala 66:30:@42386.4]
  assign _T_98696 = _T_98685[10]; // @[OneHot.scala 66:30:@42387.4]
  assign _T_98697 = _T_98685[11]; // @[OneHot.scala 66:30:@42388.4]
  assign _T_98698 = _T_98685[12]; // @[OneHot.scala 66:30:@42389.4]
  assign _T_98699 = _T_98685[13]; // @[OneHot.scala 66:30:@42390.4]
  assign _T_98700 = _T_98685[14]; // @[OneHot.scala 66:30:@42391.4]
  assign _T_98701 = _T_98685[15]; // @[OneHot.scala 66:30:@42392.4]
  assign _T_98742 = _T_97852 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42410.4]
  assign _T_98743 = _T_97849 ? 16'h4000 : _T_98742; // @[Mux.scala 31:69:@42411.4]
  assign _T_98744 = _T_97846 ? 16'h2000 : _T_98743; // @[Mux.scala 31:69:@42412.4]
  assign _T_98745 = _T_97843 ? 16'h1000 : _T_98744; // @[Mux.scala 31:69:@42413.4]
  assign _T_98746 = _T_97840 ? 16'h800 : _T_98745; // @[Mux.scala 31:69:@42414.4]
  assign _T_98747 = _T_97837 ? 16'h400 : _T_98746; // @[Mux.scala 31:69:@42415.4]
  assign _T_98748 = _T_97834 ? 16'h200 : _T_98747; // @[Mux.scala 31:69:@42416.4]
  assign _T_98749 = _T_97831 ? 16'h100 : _T_98748; // @[Mux.scala 31:69:@42417.4]
  assign _T_98750 = _T_97828 ? 16'h80 : _T_98749; // @[Mux.scala 31:69:@42418.4]
  assign _T_98751 = _T_97825 ? 16'h40 : _T_98750; // @[Mux.scala 31:69:@42419.4]
  assign _T_98752 = _T_97822 ? 16'h20 : _T_98751; // @[Mux.scala 31:69:@42420.4]
  assign _T_98753 = _T_97867 ? 16'h10 : _T_98752; // @[Mux.scala 31:69:@42421.4]
  assign _T_98754 = _T_97864 ? 16'h8 : _T_98753; // @[Mux.scala 31:69:@42422.4]
  assign _T_98755 = _T_97861 ? 16'h4 : _T_98754; // @[Mux.scala 31:69:@42423.4]
  assign _T_98756 = _T_97858 ? 16'h2 : _T_98755; // @[Mux.scala 31:69:@42424.4]
  assign _T_98757 = _T_97855 ? 16'h1 : _T_98756; // @[Mux.scala 31:69:@42425.4]
  assign _T_98758 = _T_98757[0]; // @[OneHot.scala 66:30:@42426.4]
  assign _T_98759 = _T_98757[1]; // @[OneHot.scala 66:30:@42427.4]
  assign _T_98760 = _T_98757[2]; // @[OneHot.scala 66:30:@42428.4]
  assign _T_98761 = _T_98757[3]; // @[OneHot.scala 66:30:@42429.4]
  assign _T_98762 = _T_98757[4]; // @[OneHot.scala 66:30:@42430.4]
  assign _T_98763 = _T_98757[5]; // @[OneHot.scala 66:30:@42431.4]
  assign _T_98764 = _T_98757[6]; // @[OneHot.scala 66:30:@42432.4]
  assign _T_98765 = _T_98757[7]; // @[OneHot.scala 66:30:@42433.4]
  assign _T_98766 = _T_98757[8]; // @[OneHot.scala 66:30:@42434.4]
  assign _T_98767 = _T_98757[9]; // @[OneHot.scala 66:30:@42435.4]
  assign _T_98768 = _T_98757[10]; // @[OneHot.scala 66:30:@42436.4]
  assign _T_98769 = _T_98757[11]; // @[OneHot.scala 66:30:@42437.4]
  assign _T_98770 = _T_98757[12]; // @[OneHot.scala 66:30:@42438.4]
  assign _T_98771 = _T_98757[13]; // @[OneHot.scala 66:30:@42439.4]
  assign _T_98772 = _T_98757[14]; // @[OneHot.scala 66:30:@42440.4]
  assign _T_98773 = _T_98757[15]; // @[OneHot.scala 66:30:@42441.4]
  assign _T_98814 = _T_97855 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42459.4]
  assign _T_98815 = _T_97852 ? 16'h4000 : _T_98814; // @[Mux.scala 31:69:@42460.4]
  assign _T_98816 = _T_97849 ? 16'h2000 : _T_98815; // @[Mux.scala 31:69:@42461.4]
  assign _T_98817 = _T_97846 ? 16'h1000 : _T_98816; // @[Mux.scala 31:69:@42462.4]
  assign _T_98818 = _T_97843 ? 16'h800 : _T_98817; // @[Mux.scala 31:69:@42463.4]
  assign _T_98819 = _T_97840 ? 16'h400 : _T_98818; // @[Mux.scala 31:69:@42464.4]
  assign _T_98820 = _T_97837 ? 16'h200 : _T_98819; // @[Mux.scala 31:69:@42465.4]
  assign _T_98821 = _T_97834 ? 16'h100 : _T_98820; // @[Mux.scala 31:69:@42466.4]
  assign _T_98822 = _T_97831 ? 16'h80 : _T_98821; // @[Mux.scala 31:69:@42467.4]
  assign _T_98823 = _T_97828 ? 16'h40 : _T_98822; // @[Mux.scala 31:69:@42468.4]
  assign _T_98824 = _T_97825 ? 16'h20 : _T_98823; // @[Mux.scala 31:69:@42469.4]
  assign _T_98825 = _T_97822 ? 16'h10 : _T_98824; // @[Mux.scala 31:69:@42470.4]
  assign _T_98826 = _T_97867 ? 16'h8 : _T_98825; // @[Mux.scala 31:69:@42471.4]
  assign _T_98827 = _T_97864 ? 16'h4 : _T_98826; // @[Mux.scala 31:69:@42472.4]
  assign _T_98828 = _T_97861 ? 16'h2 : _T_98827; // @[Mux.scala 31:69:@42473.4]
  assign _T_98829 = _T_97858 ? 16'h1 : _T_98828; // @[Mux.scala 31:69:@42474.4]
  assign _T_98830 = _T_98829[0]; // @[OneHot.scala 66:30:@42475.4]
  assign _T_98831 = _T_98829[1]; // @[OneHot.scala 66:30:@42476.4]
  assign _T_98832 = _T_98829[2]; // @[OneHot.scala 66:30:@42477.4]
  assign _T_98833 = _T_98829[3]; // @[OneHot.scala 66:30:@42478.4]
  assign _T_98834 = _T_98829[4]; // @[OneHot.scala 66:30:@42479.4]
  assign _T_98835 = _T_98829[5]; // @[OneHot.scala 66:30:@42480.4]
  assign _T_98836 = _T_98829[6]; // @[OneHot.scala 66:30:@42481.4]
  assign _T_98837 = _T_98829[7]; // @[OneHot.scala 66:30:@42482.4]
  assign _T_98838 = _T_98829[8]; // @[OneHot.scala 66:30:@42483.4]
  assign _T_98839 = _T_98829[9]; // @[OneHot.scala 66:30:@42484.4]
  assign _T_98840 = _T_98829[10]; // @[OneHot.scala 66:30:@42485.4]
  assign _T_98841 = _T_98829[11]; // @[OneHot.scala 66:30:@42486.4]
  assign _T_98842 = _T_98829[12]; // @[OneHot.scala 66:30:@42487.4]
  assign _T_98843 = _T_98829[13]; // @[OneHot.scala 66:30:@42488.4]
  assign _T_98844 = _T_98829[14]; // @[OneHot.scala 66:30:@42489.4]
  assign _T_98845 = _T_98829[15]; // @[OneHot.scala 66:30:@42490.4]
  assign _T_98886 = _T_97858 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42508.4]
  assign _T_98887 = _T_97855 ? 16'h4000 : _T_98886; // @[Mux.scala 31:69:@42509.4]
  assign _T_98888 = _T_97852 ? 16'h2000 : _T_98887; // @[Mux.scala 31:69:@42510.4]
  assign _T_98889 = _T_97849 ? 16'h1000 : _T_98888; // @[Mux.scala 31:69:@42511.4]
  assign _T_98890 = _T_97846 ? 16'h800 : _T_98889; // @[Mux.scala 31:69:@42512.4]
  assign _T_98891 = _T_97843 ? 16'h400 : _T_98890; // @[Mux.scala 31:69:@42513.4]
  assign _T_98892 = _T_97840 ? 16'h200 : _T_98891; // @[Mux.scala 31:69:@42514.4]
  assign _T_98893 = _T_97837 ? 16'h100 : _T_98892; // @[Mux.scala 31:69:@42515.4]
  assign _T_98894 = _T_97834 ? 16'h80 : _T_98893; // @[Mux.scala 31:69:@42516.4]
  assign _T_98895 = _T_97831 ? 16'h40 : _T_98894; // @[Mux.scala 31:69:@42517.4]
  assign _T_98896 = _T_97828 ? 16'h20 : _T_98895; // @[Mux.scala 31:69:@42518.4]
  assign _T_98897 = _T_97825 ? 16'h10 : _T_98896; // @[Mux.scala 31:69:@42519.4]
  assign _T_98898 = _T_97822 ? 16'h8 : _T_98897; // @[Mux.scala 31:69:@42520.4]
  assign _T_98899 = _T_97867 ? 16'h4 : _T_98898; // @[Mux.scala 31:69:@42521.4]
  assign _T_98900 = _T_97864 ? 16'h2 : _T_98899; // @[Mux.scala 31:69:@42522.4]
  assign _T_98901 = _T_97861 ? 16'h1 : _T_98900; // @[Mux.scala 31:69:@42523.4]
  assign _T_98902 = _T_98901[0]; // @[OneHot.scala 66:30:@42524.4]
  assign _T_98903 = _T_98901[1]; // @[OneHot.scala 66:30:@42525.4]
  assign _T_98904 = _T_98901[2]; // @[OneHot.scala 66:30:@42526.4]
  assign _T_98905 = _T_98901[3]; // @[OneHot.scala 66:30:@42527.4]
  assign _T_98906 = _T_98901[4]; // @[OneHot.scala 66:30:@42528.4]
  assign _T_98907 = _T_98901[5]; // @[OneHot.scala 66:30:@42529.4]
  assign _T_98908 = _T_98901[6]; // @[OneHot.scala 66:30:@42530.4]
  assign _T_98909 = _T_98901[7]; // @[OneHot.scala 66:30:@42531.4]
  assign _T_98910 = _T_98901[8]; // @[OneHot.scala 66:30:@42532.4]
  assign _T_98911 = _T_98901[9]; // @[OneHot.scala 66:30:@42533.4]
  assign _T_98912 = _T_98901[10]; // @[OneHot.scala 66:30:@42534.4]
  assign _T_98913 = _T_98901[11]; // @[OneHot.scala 66:30:@42535.4]
  assign _T_98914 = _T_98901[12]; // @[OneHot.scala 66:30:@42536.4]
  assign _T_98915 = _T_98901[13]; // @[OneHot.scala 66:30:@42537.4]
  assign _T_98916 = _T_98901[14]; // @[OneHot.scala 66:30:@42538.4]
  assign _T_98917 = _T_98901[15]; // @[OneHot.scala 66:30:@42539.4]
  assign _T_98958 = _T_97861 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42557.4]
  assign _T_98959 = _T_97858 ? 16'h4000 : _T_98958; // @[Mux.scala 31:69:@42558.4]
  assign _T_98960 = _T_97855 ? 16'h2000 : _T_98959; // @[Mux.scala 31:69:@42559.4]
  assign _T_98961 = _T_97852 ? 16'h1000 : _T_98960; // @[Mux.scala 31:69:@42560.4]
  assign _T_98962 = _T_97849 ? 16'h800 : _T_98961; // @[Mux.scala 31:69:@42561.4]
  assign _T_98963 = _T_97846 ? 16'h400 : _T_98962; // @[Mux.scala 31:69:@42562.4]
  assign _T_98964 = _T_97843 ? 16'h200 : _T_98963; // @[Mux.scala 31:69:@42563.4]
  assign _T_98965 = _T_97840 ? 16'h100 : _T_98964; // @[Mux.scala 31:69:@42564.4]
  assign _T_98966 = _T_97837 ? 16'h80 : _T_98965; // @[Mux.scala 31:69:@42565.4]
  assign _T_98967 = _T_97834 ? 16'h40 : _T_98966; // @[Mux.scala 31:69:@42566.4]
  assign _T_98968 = _T_97831 ? 16'h20 : _T_98967; // @[Mux.scala 31:69:@42567.4]
  assign _T_98969 = _T_97828 ? 16'h10 : _T_98968; // @[Mux.scala 31:69:@42568.4]
  assign _T_98970 = _T_97825 ? 16'h8 : _T_98969; // @[Mux.scala 31:69:@42569.4]
  assign _T_98971 = _T_97822 ? 16'h4 : _T_98970; // @[Mux.scala 31:69:@42570.4]
  assign _T_98972 = _T_97867 ? 16'h2 : _T_98971; // @[Mux.scala 31:69:@42571.4]
  assign _T_98973 = _T_97864 ? 16'h1 : _T_98972; // @[Mux.scala 31:69:@42572.4]
  assign _T_98974 = _T_98973[0]; // @[OneHot.scala 66:30:@42573.4]
  assign _T_98975 = _T_98973[1]; // @[OneHot.scala 66:30:@42574.4]
  assign _T_98976 = _T_98973[2]; // @[OneHot.scala 66:30:@42575.4]
  assign _T_98977 = _T_98973[3]; // @[OneHot.scala 66:30:@42576.4]
  assign _T_98978 = _T_98973[4]; // @[OneHot.scala 66:30:@42577.4]
  assign _T_98979 = _T_98973[5]; // @[OneHot.scala 66:30:@42578.4]
  assign _T_98980 = _T_98973[6]; // @[OneHot.scala 66:30:@42579.4]
  assign _T_98981 = _T_98973[7]; // @[OneHot.scala 66:30:@42580.4]
  assign _T_98982 = _T_98973[8]; // @[OneHot.scala 66:30:@42581.4]
  assign _T_98983 = _T_98973[9]; // @[OneHot.scala 66:30:@42582.4]
  assign _T_98984 = _T_98973[10]; // @[OneHot.scala 66:30:@42583.4]
  assign _T_98985 = _T_98973[11]; // @[OneHot.scala 66:30:@42584.4]
  assign _T_98986 = _T_98973[12]; // @[OneHot.scala 66:30:@42585.4]
  assign _T_98987 = _T_98973[13]; // @[OneHot.scala 66:30:@42586.4]
  assign _T_98988 = _T_98973[14]; // @[OneHot.scala 66:30:@42587.4]
  assign _T_98989 = _T_98973[15]; // @[OneHot.scala 66:30:@42588.4]
  assign _T_99030 = _T_97864 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42606.4]
  assign _T_99031 = _T_97861 ? 16'h4000 : _T_99030; // @[Mux.scala 31:69:@42607.4]
  assign _T_99032 = _T_97858 ? 16'h2000 : _T_99031; // @[Mux.scala 31:69:@42608.4]
  assign _T_99033 = _T_97855 ? 16'h1000 : _T_99032; // @[Mux.scala 31:69:@42609.4]
  assign _T_99034 = _T_97852 ? 16'h800 : _T_99033; // @[Mux.scala 31:69:@42610.4]
  assign _T_99035 = _T_97849 ? 16'h400 : _T_99034; // @[Mux.scala 31:69:@42611.4]
  assign _T_99036 = _T_97846 ? 16'h200 : _T_99035; // @[Mux.scala 31:69:@42612.4]
  assign _T_99037 = _T_97843 ? 16'h100 : _T_99036; // @[Mux.scala 31:69:@42613.4]
  assign _T_99038 = _T_97840 ? 16'h80 : _T_99037; // @[Mux.scala 31:69:@42614.4]
  assign _T_99039 = _T_97837 ? 16'h40 : _T_99038; // @[Mux.scala 31:69:@42615.4]
  assign _T_99040 = _T_97834 ? 16'h20 : _T_99039; // @[Mux.scala 31:69:@42616.4]
  assign _T_99041 = _T_97831 ? 16'h10 : _T_99040; // @[Mux.scala 31:69:@42617.4]
  assign _T_99042 = _T_97828 ? 16'h8 : _T_99041; // @[Mux.scala 31:69:@42618.4]
  assign _T_99043 = _T_97825 ? 16'h4 : _T_99042; // @[Mux.scala 31:69:@42619.4]
  assign _T_99044 = _T_97822 ? 16'h2 : _T_99043; // @[Mux.scala 31:69:@42620.4]
  assign _T_99045 = _T_97867 ? 16'h1 : _T_99044; // @[Mux.scala 31:69:@42621.4]
  assign _T_99046 = _T_99045[0]; // @[OneHot.scala 66:30:@42622.4]
  assign _T_99047 = _T_99045[1]; // @[OneHot.scala 66:30:@42623.4]
  assign _T_99048 = _T_99045[2]; // @[OneHot.scala 66:30:@42624.4]
  assign _T_99049 = _T_99045[3]; // @[OneHot.scala 66:30:@42625.4]
  assign _T_99050 = _T_99045[4]; // @[OneHot.scala 66:30:@42626.4]
  assign _T_99051 = _T_99045[5]; // @[OneHot.scala 66:30:@42627.4]
  assign _T_99052 = _T_99045[6]; // @[OneHot.scala 66:30:@42628.4]
  assign _T_99053 = _T_99045[7]; // @[OneHot.scala 66:30:@42629.4]
  assign _T_99054 = _T_99045[8]; // @[OneHot.scala 66:30:@42630.4]
  assign _T_99055 = _T_99045[9]; // @[OneHot.scala 66:30:@42631.4]
  assign _T_99056 = _T_99045[10]; // @[OneHot.scala 66:30:@42632.4]
  assign _T_99057 = _T_99045[11]; // @[OneHot.scala 66:30:@42633.4]
  assign _T_99058 = _T_99045[12]; // @[OneHot.scala 66:30:@42634.4]
  assign _T_99059 = _T_99045[13]; // @[OneHot.scala 66:30:@42635.4]
  assign _T_99060 = _T_99045[14]; // @[OneHot.scala 66:30:@42636.4]
  assign _T_99061 = _T_99045[15]; // @[OneHot.scala 66:30:@42637.4]
  assign _T_99126 = {_T_97973,_T_97972,_T_97971,_T_97970,_T_97969,_T_97968,_T_97967,_T_97966}; // @[Mux.scala 19:72:@42661.4]
  assign _T_99134 = {_T_97981,_T_97980,_T_97979,_T_97978,_T_97977,_T_97976,_T_97975,_T_97974,_T_99126}; // @[Mux.scala 19:72:@42669.4]
  assign _T_99136 = _T_90408 ? _T_99134 : 16'h0; // @[Mux.scala 19:72:@42670.4]
  assign _T_99143 = {_T_98044,_T_98043,_T_98042,_T_98041,_T_98040,_T_98039,_T_98038,_T_98053}; // @[Mux.scala 19:72:@42677.4]
  assign _T_99151 = {_T_98052,_T_98051,_T_98050,_T_98049,_T_98048,_T_98047,_T_98046,_T_98045,_T_99143}; // @[Mux.scala 19:72:@42685.4]
  assign _T_99153 = _T_90409 ? _T_99151 : 16'h0; // @[Mux.scala 19:72:@42686.4]
  assign _T_99160 = {_T_98115,_T_98114,_T_98113,_T_98112,_T_98111,_T_98110,_T_98125,_T_98124}; // @[Mux.scala 19:72:@42693.4]
  assign _T_99168 = {_T_98123,_T_98122,_T_98121,_T_98120,_T_98119,_T_98118,_T_98117,_T_98116,_T_99160}; // @[Mux.scala 19:72:@42701.4]
  assign _T_99170 = _T_90410 ? _T_99168 : 16'h0; // @[Mux.scala 19:72:@42702.4]
  assign _T_99177 = {_T_98186,_T_98185,_T_98184,_T_98183,_T_98182,_T_98197,_T_98196,_T_98195}; // @[Mux.scala 19:72:@42709.4]
  assign _T_99185 = {_T_98194,_T_98193,_T_98192,_T_98191,_T_98190,_T_98189,_T_98188,_T_98187,_T_99177}; // @[Mux.scala 19:72:@42717.4]
  assign _T_99187 = _T_90411 ? _T_99185 : 16'h0; // @[Mux.scala 19:72:@42718.4]
  assign _T_99194 = {_T_98257,_T_98256,_T_98255,_T_98254,_T_98269,_T_98268,_T_98267,_T_98266}; // @[Mux.scala 19:72:@42725.4]
  assign _T_99202 = {_T_98265,_T_98264,_T_98263,_T_98262,_T_98261,_T_98260,_T_98259,_T_98258,_T_99194}; // @[Mux.scala 19:72:@42733.4]
  assign _T_99204 = _T_90412 ? _T_99202 : 16'h0; // @[Mux.scala 19:72:@42734.4]
  assign _T_99211 = {_T_98328,_T_98327,_T_98326,_T_98341,_T_98340,_T_98339,_T_98338,_T_98337}; // @[Mux.scala 19:72:@42741.4]
  assign _T_99219 = {_T_98336,_T_98335,_T_98334,_T_98333,_T_98332,_T_98331,_T_98330,_T_98329,_T_99211}; // @[Mux.scala 19:72:@42749.4]
  assign _T_99221 = _T_90413 ? _T_99219 : 16'h0; // @[Mux.scala 19:72:@42750.4]
  assign _T_99228 = {_T_98399,_T_98398,_T_98413,_T_98412,_T_98411,_T_98410,_T_98409,_T_98408}; // @[Mux.scala 19:72:@42757.4]
  assign _T_99236 = {_T_98407,_T_98406,_T_98405,_T_98404,_T_98403,_T_98402,_T_98401,_T_98400,_T_99228}; // @[Mux.scala 19:72:@42765.4]
  assign _T_99238 = _T_90414 ? _T_99236 : 16'h0; // @[Mux.scala 19:72:@42766.4]
  assign _T_99245 = {_T_98470,_T_98485,_T_98484,_T_98483,_T_98482,_T_98481,_T_98480,_T_98479}; // @[Mux.scala 19:72:@42773.4]
  assign _T_99253 = {_T_98478,_T_98477,_T_98476,_T_98475,_T_98474,_T_98473,_T_98472,_T_98471,_T_99245}; // @[Mux.scala 19:72:@42781.4]
  assign _T_99255 = _T_90415 ? _T_99253 : 16'h0; // @[Mux.scala 19:72:@42782.4]
  assign _T_99262 = {_T_98557,_T_98556,_T_98555,_T_98554,_T_98553,_T_98552,_T_98551,_T_98550}; // @[Mux.scala 19:72:@42789.4]
  assign _T_99270 = {_T_98549,_T_98548,_T_98547,_T_98546,_T_98545,_T_98544,_T_98543,_T_98542,_T_99262}; // @[Mux.scala 19:72:@42797.4]
  assign _T_99272 = _T_90416 ? _T_99270 : 16'h0; // @[Mux.scala 19:72:@42798.4]
  assign _T_99279 = {_T_98628,_T_98627,_T_98626,_T_98625,_T_98624,_T_98623,_T_98622,_T_98621}; // @[Mux.scala 19:72:@42805.4]
  assign _T_99287 = {_T_98620,_T_98619,_T_98618,_T_98617,_T_98616,_T_98615,_T_98614,_T_98629,_T_99279}; // @[Mux.scala 19:72:@42813.4]
  assign _T_99289 = _T_90417 ? _T_99287 : 16'h0; // @[Mux.scala 19:72:@42814.4]
  assign _T_99296 = {_T_98699,_T_98698,_T_98697,_T_98696,_T_98695,_T_98694,_T_98693,_T_98692}; // @[Mux.scala 19:72:@42821.4]
  assign _T_99304 = {_T_98691,_T_98690,_T_98689,_T_98688,_T_98687,_T_98686,_T_98701,_T_98700,_T_99296}; // @[Mux.scala 19:72:@42829.4]
  assign _T_99306 = _T_90418 ? _T_99304 : 16'h0; // @[Mux.scala 19:72:@42830.4]
  assign _T_99313 = {_T_98770,_T_98769,_T_98768,_T_98767,_T_98766,_T_98765,_T_98764,_T_98763}; // @[Mux.scala 19:72:@42837.4]
  assign _T_99321 = {_T_98762,_T_98761,_T_98760,_T_98759,_T_98758,_T_98773,_T_98772,_T_98771,_T_99313}; // @[Mux.scala 19:72:@42845.4]
  assign _T_99323 = _T_90419 ? _T_99321 : 16'h0; // @[Mux.scala 19:72:@42846.4]
  assign _T_99330 = {_T_98841,_T_98840,_T_98839,_T_98838,_T_98837,_T_98836,_T_98835,_T_98834}; // @[Mux.scala 19:72:@42853.4]
  assign _T_99338 = {_T_98833,_T_98832,_T_98831,_T_98830,_T_98845,_T_98844,_T_98843,_T_98842,_T_99330}; // @[Mux.scala 19:72:@42861.4]
  assign _T_99340 = _T_90420 ? _T_99338 : 16'h0; // @[Mux.scala 19:72:@42862.4]
  assign _T_99347 = {_T_98912,_T_98911,_T_98910,_T_98909,_T_98908,_T_98907,_T_98906,_T_98905}; // @[Mux.scala 19:72:@42869.4]
  assign _T_99355 = {_T_98904,_T_98903,_T_98902,_T_98917,_T_98916,_T_98915,_T_98914,_T_98913,_T_99347}; // @[Mux.scala 19:72:@42877.4]
  assign _T_99357 = _T_90421 ? _T_99355 : 16'h0; // @[Mux.scala 19:72:@42878.4]
  assign _T_99364 = {_T_98983,_T_98982,_T_98981,_T_98980,_T_98979,_T_98978,_T_98977,_T_98976}; // @[Mux.scala 19:72:@42885.4]
  assign _T_99372 = {_T_98975,_T_98974,_T_98989,_T_98988,_T_98987,_T_98986,_T_98985,_T_98984,_T_99364}; // @[Mux.scala 19:72:@42893.4]
  assign _T_99374 = _T_90422 ? _T_99372 : 16'h0; // @[Mux.scala 19:72:@42894.4]
  assign _T_99381 = {_T_99054,_T_99053,_T_99052,_T_99051,_T_99050,_T_99049,_T_99048,_T_99047}; // @[Mux.scala 19:72:@42901.4]
  assign _T_99389 = {_T_99046,_T_99061,_T_99060,_T_99059,_T_99058,_T_99057,_T_99056,_T_99055,_T_99381}; // @[Mux.scala 19:72:@42909.4]
  assign _T_99391 = _T_90423 ? _T_99389 : 16'h0; // @[Mux.scala 19:72:@42910.4]
  assign _T_99392 = _T_99136 | _T_99153; // @[Mux.scala 19:72:@42911.4]
  assign _T_99393 = _T_99392 | _T_99170; // @[Mux.scala 19:72:@42912.4]
  assign _T_99394 = _T_99393 | _T_99187; // @[Mux.scala 19:72:@42913.4]
  assign _T_99395 = _T_99394 | _T_99204; // @[Mux.scala 19:72:@42914.4]
  assign _T_99396 = _T_99395 | _T_99221; // @[Mux.scala 19:72:@42915.4]
  assign _T_99397 = _T_99396 | _T_99238; // @[Mux.scala 19:72:@42916.4]
  assign _T_99398 = _T_99397 | _T_99255; // @[Mux.scala 19:72:@42917.4]
  assign _T_99399 = _T_99398 | _T_99272; // @[Mux.scala 19:72:@42918.4]
  assign _T_99400 = _T_99399 | _T_99289; // @[Mux.scala 19:72:@42919.4]
  assign _T_99401 = _T_99400 | _T_99306; // @[Mux.scala 19:72:@42920.4]
  assign _T_99402 = _T_99401 | _T_99323; // @[Mux.scala 19:72:@42921.4]
  assign _T_99403 = _T_99402 | _T_99340; // @[Mux.scala 19:72:@42922.4]
  assign _T_99404 = _T_99403 | _T_99357; // @[Mux.scala 19:72:@42923.4]
  assign _T_99405 = _T_99404 | _T_99374; // @[Mux.scala 19:72:@42924.4]
  assign _T_99406 = _T_99405 | _T_99391; // @[Mux.scala 19:72:@42925.4]
  assign inputPriorityPorts_1_0 = _T_99406[0]; // @[Mux.scala 19:72:@42929.4]
  assign inputPriorityPorts_1_1 = _T_99406[1]; // @[Mux.scala 19:72:@42931.4]
  assign inputPriorityPorts_1_2 = _T_99406[2]; // @[Mux.scala 19:72:@42933.4]
  assign inputPriorityPorts_1_3 = _T_99406[3]; // @[Mux.scala 19:72:@42935.4]
  assign inputPriorityPorts_1_4 = _T_99406[4]; // @[Mux.scala 19:72:@42937.4]
  assign inputPriorityPorts_1_5 = _T_99406[5]; // @[Mux.scala 19:72:@42939.4]
  assign inputPriorityPorts_1_6 = _T_99406[6]; // @[Mux.scala 19:72:@42941.4]
  assign inputPriorityPorts_1_7 = _T_99406[7]; // @[Mux.scala 19:72:@42943.4]
  assign inputPriorityPorts_1_8 = _T_99406[8]; // @[Mux.scala 19:72:@42945.4]
  assign inputPriorityPorts_1_9 = _T_99406[9]; // @[Mux.scala 19:72:@42947.4]
  assign inputPriorityPorts_1_10 = _T_99406[10]; // @[Mux.scala 19:72:@42949.4]
  assign inputPriorityPorts_1_11 = _T_99406[11]; // @[Mux.scala 19:72:@42951.4]
  assign inputPriorityPorts_1_12 = _T_99406[12]; // @[Mux.scala 19:72:@42953.4]
  assign inputPriorityPorts_1_13 = _T_99406[13]; // @[Mux.scala 19:72:@42955.4]
  assign inputPriorityPorts_1_14 = _T_99406[14]; // @[Mux.scala 19:72:@42957.4]
  assign inputPriorityPorts_1_15 = _T_99406[15]; // @[Mux.scala 19:72:@42959.4]
  assign _T_99608 = portQ_15 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43013.4]
  assign _T_99609 = portQ_14 ? 16'h4000 : _T_99608; // @[Mux.scala 31:69:@43014.4]
  assign _T_99610 = portQ_13 ? 16'h2000 : _T_99609; // @[Mux.scala 31:69:@43015.4]
  assign _T_99611 = portQ_12 ? 16'h1000 : _T_99610; // @[Mux.scala 31:69:@43016.4]
  assign _T_99612 = portQ_11 ? 16'h800 : _T_99611; // @[Mux.scala 31:69:@43017.4]
  assign _T_99613 = portQ_10 ? 16'h400 : _T_99612; // @[Mux.scala 31:69:@43018.4]
  assign _T_99614 = portQ_9 ? 16'h200 : _T_99613; // @[Mux.scala 31:69:@43019.4]
  assign _T_99615 = portQ_8 ? 16'h100 : _T_99614; // @[Mux.scala 31:69:@43020.4]
  assign _T_99616 = portQ_7 ? 16'h80 : _T_99615; // @[Mux.scala 31:69:@43021.4]
  assign _T_99617 = portQ_6 ? 16'h40 : _T_99616; // @[Mux.scala 31:69:@43022.4]
  assign _T_99618 = portQ_5 ? 16'h20 : _T_99617; // @[Mux.scala 31:69:@43023.4]
  assign _T_99619 = portQ_4 ? 16'h10 : _T_99618; // @[Mux.scala 31:69:@43024.4]
  assign _T_99620 = portQ_3 ? 16'h8 : _T_99619; // @[Mux.scala 31:69:@43025.4]
  assign _T_99621 = portQ_2 ? 16'h4 : _T_99620; // @[Mux.scala 31:69:@43026.4]
  assign _T_99622 = portQ_1 ? 16'h2 : _T_99621; // @[Mux.scala 31:69:@43027.4]
  assign _T_99623 = portQ_0 ? 16'h1 : _T_99622; // @[Mux.scala 31:69:@43028.4]
  assign _T_99624 = _T_99623[0]; // @[OneHot.scala 66:30:@43029.4]
  assign _T_99625 = _T_99623[1]; // @[OneHot.scala 66:30:@43030.4]
  assign _T_99626 = _T_99623[2]; // @[OneHot.scala 66:30:@43031.4]
  assign _T_99627 = _T_99623[3]; // @[OneHot.scala 66:30:@43032.4]
  assign _T_99628 = _T_99623[4]; // @[OneHot.scala 66:30:@43033.4]
  assign _T_99629 = _T_99623[5]; // @[OneHot.scala 66:30:@43034.4]
  assign _T_99630 = _T_99623[6]; // @[OneHot.scala 66:30:@43035.4]
  assign _T_99631 = _T_99623[7]; // @[OneHot.scala 66:30:@43036.4]
  assign _T_99632 = _T_99623[8]; // @[OneHot.scala 66:30:@43037.4]
  assign _T_99633 = _T_99623[9]; // @[OneHot.scala 66:30:@43038.4]
  assign _T_99634 = _T_99623[10]; // @[OneHot.scala 66:30:@43039.4]
  assign _T_99635 = _T_99623[11]; // @[OneHot.scala 66:30:@43040.4]
  assign _T_99636 = _T_99623[12]; // @[OneHot.scala 66:30:@43041.4]
  assign _T_99637 = _T_99623[13]; // @[OneHot.scala 66:30:@43042.4]
  assign _T_99638 = _T_99623[14]; // @[OneHot.scala 66:30:@43043.4]
  assign _T_99639 = _T_99623[15]; // @[OneHot.scala 66:30:@43044.4]
  assign _T_99680 = portQ_0 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43062.4]
  assign _T_99681 = portQ_15 ? 16'h4000 : _T_99680; // @[Mux.scala 31:69:@43063.4]
  assign _T_99682 = portQ_14 ? 16'h2000 : _T_99681; // @[Mux.scala 31:69:@43064.4]
  assign _T_99683 = portQ_13 ? 16'h1000 : _T_99682; // @[Mux.scala 31:69:@43065.4]
  assign _T_99684 = portQ_12 ? 16'h800 : _T_99683; // @[Mux.scala 31:69:@43066.4]
  assign _T_99685 = portQ_11 ? 16'h400 : _T_99684; // @[Mux.scala 31:69:@43067.4]
  assign _T_99686 = portQ_10 ? 16'h200 : _T_99685; // @[Mux.scala 31:69:@43068.4]
  assign _T_99687 = portQ_9 ? 16'h100 : _T_99686; // @[Mux.scala 31:69:@43069.4]
  assign _T_99688 = portQ_8 ? 16'h80 : _T_99687; // @[Mux.scala 31:69:@43070.4]
  assign _T_99689 = portQ_7 ? 16'h40 : _T_99688; // @[Mux.scala 31:69:@43071.4]
  assign _T_99690 = portQ_6 ? 16'h20 : _T_99689; // @[Mux.scala 31:69:@43072.4]
  assign _T_99691 = portQ_5 ? 16'h10 : _T_99690; // @[Mux.scala 31:69:@43073.4]
  assign _T_99692 = portQ_4 ? 16'h8 : _T_99691; // @[Mux.scala 31:69:@43074.4]
  assign _T_99693 = portQ_3 ? 16'h4 : _T_99692; // @[Mux.scala 31:69:@43075.4]
  assign _T_99694 = portQ_2 ? 16'h2 : _T_99693; // @[Mux.scala 31:69:@43076.4]
  assign _T_99695 = portQ_1 ? 16'h1 : _T_99694; // @[Mux.scala 31:69:@43077.4]
  assign _T_99696 = _T_99695[0]; // @[OneHot.scala 66:30:@43078.4]
  assign _T_99697 = _T_99695[1]; // @[OneHot.scala 66:30:@43079.4]
  assign _T_99698 = _T_99695[2]; // @[OneHot.scala 66:30:@43080.4]
  assign _T_99699 = _T_99695[3]; // @[OneHot.scala 66:30:@43081.4]
  assign _T_99700 = _T_99695[4]; // @[OneHot.scala 66:30:@43082.4]
  assign _T_99701 = _T_99695[5]; // @[OneHot.scala 66:30:@43083.4]
  assign _T_99702 = _T_99695[6]; // @[OneHot.scala 66:30:@43084.4]
  assign _T_99703 = _T_99695[7]; // @[OneHot.scala 66:30:@43085.4]
  assign _T_99704 = _T_99695[8]; // @[OneHot.scala 66:30:@43086.4]
  assign _T_99705 = _T_99695[9]; // @[OneHot.scala 66:30:@43087.4]
  assign _T_99706 = _T_99695[10]; // @[OneHot.scala 66:30:@43088.4]
  assign _T_99707 = _T_99695[11]; // @[OneHot.scala 66:30:@43089.4]
  assign _T_99708 = _T_99695[12]; // @[OneHot.scala 66:30:@43090.4]
  assign _T_99709 = _T_99695[13]; // @[OneHot.scala 66:30:@43091.4]
  assign _T_99710 = _T_99695[14]; // @[OneHot.scala 66:30:@43092.4]
  assign _T_99711 = _T_99695[15]; // @[OneHot.scala 66:30:@43093.4]
  assign _T_99752 = portQ_1 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43111.4]
  assign _T_99753 = portQ_0 ? 16'h4000 : _T_99752; // @[Mux.scala 31:69:@43112.4]
  assign _T_99754 = portQ_15 ? 16'h2000 : _T_99753; // @[Mux.scala 31:69:@43113.4]
  assign _T_99755 = portQ_14 ? 16'h1000 : _T_99754; // @[Mux.scala 31:69:@43114.4]
  assign _T_99756 = portQ_13 ? 16'h800 : _T_99755; // @[Mux.scala 31:69:@43115.4]
  assign _T_99757 = portQ_12 ? 16'h400 : _T_99756; // @[Mux.scala 31:69:@43116.4]
  assign _T_99758 = portQ_11 ? 16'h200 : _T_99757; // @[Mux.scala 31:69:@43117.4]
  assign _T_99759 = portQ_10 ? 16'h100 : _T_99758; // @[Mux.scala 31:69:@43118.4]
  assign _T_99760 = portQ_9 ? 16'h80 : _T_99759; // @[Mux.scala 31:69:@43119.4]
  assign _T_99761 = portQ_8 ? 16'h40 : _T_99760; // @[Mux.scala 31:69:@43120.4]
  assign _T_99762 = portQ_7 ? 16'h20 : _T_99761; // @[Mux.scala 31:69:@43121.4]
  assign _T_99763 = portQ_6 ? 16'h10 : _T_99762; // @[Mux.scala 31:69:@43122.4]
  assign _T_99764 = portQ_5 ? 16'h8 : _T_99763; // @[Mux.scala 31:69:@43123.4]
  assign _T_99765 = portQ_4 ? 16'h4 : _T_99764; // @[Mux.scala 31:69:@43124.4]
  assign _T_99766 = portQ_3 ? 16'h2 : _T_99765; // @[Mux.scala 31:69:@43125.4]
  assign _T_99767 = portQ_2 ? 16'h1 : _T_99766; // @[Mux.scala 31:69:@43126.4]
  assign _T_99768 = _T_99767[0]; // @[OneHot.scala 66:30:@43127.4]
  assign _T_99769 = _T_99767[1]; // @[OneHot.scala 66:30:@43128.4]
  assign _T_99770 = _T_99767[2]; // @[OneHot.scala 66:30:@43129.4]
  assign _T_99771 = _T_99767[3]; // @[OneHot.scala 66:30:@43130.4]
  assign _T_99772 = _T_99767[4]; // @[OneHot.scala 66:30:@43131.4]
  assign _T_99773 = _T_99767[5]; // @[OneHot.scala 66:30:@43132.4]
  assign _T_99774 = _T_99767[6]; // @[OneHot.scala 66:30:@43133.4]
  assign _T_99775 = _T_99767[7]; // @[OneHot.scala 66:30:@43134.4]
  assign _T_99776 = _T_99767[8]; // @[OneHot.scala 66:30:@43135.4]
  assign _T_99777 = _T_99767[9]; // @[OneHot.scala 66:30:@43136.4]
  assign _T_99778 = _T_99767[10]; // @[OneHot.scala 66:30:@43137.4]
  assign _T_99779 = _T_99767[11]; // @[OneHot.scala 66:30:@43138.4]
  assign _T_99780 = _T_99767[12]; // @[OneHot.scala 66:30:@43139.4]
  assign _T_99781 = _T_99767[13]; // @[OneHot.scala 66:30:@43140.4]
  assign _T_99782 = _T_99767[14]; // @[OneHot.scala 66:30:@43141.4]
  assign _T_99783 = _T_99767[15]; // @[OneHot.scala 66:30:@43142.4]
  assign _T_99824 = portQ_2 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43160.4]
  assign _T_99825 = portQ_1 ? 16'h4000 : _T_99824; // @[Mux.scala 31:69:@43161.4]
  assign _T_99826 = portQ_0 ? 16'h2000 : _T_99825; // @[Mux.scala 31:69:@43162.4]
  assign _T_99827 = portQ_15 ? 16'h1000 : _T_99826; // @[Mux.scala 31:69:@43163.4]
  assign _T_99828 = portQ_14 ? 16'h800 : _T_99827; // @[Mux.scala 31:69:@43164.4]
  assign _T_99829 = portQ_13 ? 16'h400 : _T_99828; // @[Mux.scala 31:69:@43165.4]
  assign _T_99830 = portQ_12 ? 16'h200 : _T_99829; // @[Mux.scala 31:69:@43166.4]
  assign _T_99831 = portQ_11 ? 16'h100 : _T_99830; // @[Mux.scala 31:69:@43167.4]
  assign _T_99832 = portQ_10 ? 16'h80 : _T_99831; // @[Mux.scala 31:69:@43168.4]
  assign _T_99833 = portQ_9 ? 16'h40 : _T_99832; // @[Mux.scala 31:69:@43169.4]
  assign _T_99834 = portQ_8 ? 16'h20 : _T_99833; // @[Mux.scala 31:69:@43170.4]
  assign _T_99835 = portQ_7 ? 16'h10 : _T_99834; // @[Mux.scala 31:69:@43171.4]
  assign _T_99836 = portQ_6 ? 16'h8 : _T_99835; // @[Mux.scala 31:69:@43172.4]
  assign _T_99837 = portQ_5 ? 16'h4 : _T_99836; // @[Mux.scala 31:69:@43173.4]
  assign _T_99838 = portQ_4 ? 16'h2 : _T_99837; // @[Mux.scala 31:69:@43174.4]
  assign _T_99839 = portQ_3 ? 16'h1 : _T_99838; // @[Mux.scala 31:69:@43175.4]
  assign _T_99840 = _T_99839[0]; // @[OneHot.scala 66:30:@43176.4]
  assign _T_99841 = _T_99839[1]; // @[OneHot.scala 66:30:@43177.4]
  assign _T_99842 = _T_99839[2]; // @[OneHot.scala 66:30:@43178.4]
  assign _T_99843 = _T_99839[3]; // @[OneHot.scala 66:30:@43179.4]
  assign _T_99844 = _T_99839[4]; // @[OneHot.scala 66:30:@43180.4]
  assign _T_99845 = _T_99839[5]; // @[OneHot.scala 66:30:@43181.4]
  assign _T_99846 = _T_99839[6]; // @[OneHot.scala 66:30:@43182.4]
  assign _T_99847 = _T_99839[7]; // @[OneHot.scala 66:30:@43183.4]
  assign _T_99848 = _T_99839[8]; // @[OneHot.scala 66:30:@43184.4]
  assign _T_99849 = _T_99839[9]; // @[OneHot.scala 66:30:@43185.4]
  assign _T_99850 = _T_99839[10]; // @[OneHot.scala 66:30:@43186.4]
  assign _T_99851 = _T_99839[11]; // @[OneHot.scala 66:30:@43187.4]
  assign _T_99852 = _T_99839[12]; // @[OneHot.scala 66:30:@43188.4]
  assign _T_99853 = _T_99839[13]; // @[OneHot.scala 66:30:@43189.4]
  assign _T_99854 = _T_99839[14]; // @[OneHot.scala 66:30:@43190.4]
  assign _T_99855 = _T_99839[15]; // @[OneHot.scala 66:30:@43191.4]
  assign _T_99896 = portQ_3 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43209.4]
  assign _T_99897 = portQ_2 ? 16'h4000 : _T_99896; // @[Mux.scala 31:69:@43210.4]
  assign _T_99898 = portQ_1 ? 16'h2000 : _T_99897; // @[Mux.scala 31:69:@43211.4]
  assign _T_99899 = portQ_0 ? 16'h1000 : _T_99898; // @[Mux.scala 31:69:@43212.4]
  assign _T_99900 = portQ_15 ? 16'h800 : _T_99899; // @[Mux.scala 31:69:@43213.4]
  assign _T_99901 = portQ_14 ? 16'h400 : _T_99900; // @[Mux.scala 31:69:@43214.4]
  assign _T_99902 = portQ_13 ? 16'h200 : _T_99901; // @[Mux.scala 31:69:@43215.4]
  assign _T_99903 = portQ_12 ? 16'h100 : _T_99902; // @[Mux.scala 31:69:@43216.4]
  assign _T_99904 = portQ_11 ? 16'h80 : _T_99903; // @[Mux.scala 31:69:@43217.4]
  assign _T_99905 = portQ_10 ? 16'h40 : _T_99904; // @[Mux.scala 31:69:@43218.4]
  assign _T_99906 = portQ_9 ? 16'h20 : _T_99905; // @[Mux.scala 31:69:@43219.4]
  assign _T_99907 = portQ_8 ? 16'h10 : _T_99906; // @[Mux.scala 31:69:@43220.4]
  assign _T_99908 = portQ_7 ? 16'h8 : _T_99907; // @[Mux.scala 31:69:@43221.4]
  assign _T_99909 = portQ_6 ? 16'h4 : _T_99908; // @[Mux.scala 31:69:@43222.4]
  assign _T_99910 = portQ_5 ? 16'h2 : _T_99909; // @[Mux.scala 31:69:@43223.4]
  assign _T_99911 = portQ_4 ? 16'h1 : _T_99910; // @[Mux.scala 31:69:@43224.4]
  assign _T_99912 = _T_99911[0]; // @[OneHot.scala 66:30:@43225.4]
  assign _T_99913 = _T_99911[1]; // @[OneHot.scala 66:30:@43226.4]
  assign _T_99914 = _T_99911[2]; // @[OneHot.scala 66:30:@43227.4]
  assign _T_99915 = _T_99911[3]; // @[OneHot.scala 66:30:@43228.4]
  assign _T_99916 = _T_99911[4]; // @[OneHot.scala 66:30:@43229.4]
  assign _T_99917 = _T_99911[5]; // @[OneHot.scala 66:30:@43230.4]
  assign _T_99918 = _T_99911[6]; // @[OneHot.scala 66:30:@43231.4]
  assign _T_99919 = _T_99911[7]; // @[OneHot.scala 66:30:@43232.4]
  assign _T_99920 = _T_99911[8]; // @[OneHot.scala 66:30:@43233.4]
  assign _T_99921 = _T_99911[9]; // @[OneHot.scala 66:30:@43234.4]
  assign _T_99922 = _T_99911[10]; // @[OneHot.scala 66:30:@43235.4]
  assign _T_99923 = _T_99911[11]; // @[OneHot.scala 66:30:@43236.4]
  assign _T_99924 = _T_99911[12]; // @[OneHot.scala 66:30:@43237.4]
  assign _T_99925 = _T_99911[13]; // @[OneHot.scala 66:30:@43238.4]
  assign _T_99926 = _T_99911[14]; // @[OneHot.scala 66:30:@43239.4]
  assign _T_99927 = _T_99911[15]; // @[OneHot.scala 66:30:@43240.4]
  assign _T_99968 = portQ_4 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43258.4]
  assign _T_99969 = portQ_3 ? 16'h4000 : _T_99968; // @[Mux.scala 31:69:@43259.4]
  assign _T_99970 = portQ_2 ? 16'h2000 : _T_99969; // @[Mux.scala 31:69:@43260.4]
  assign _T_99971 = portQ_1 ? 16'h1000 : _T_99970; // @[Mux.scala 31:69:@43261.4]
  assign _T_99972 = portQ_0 ? 16'h800 : _T_99971; // @[Mux.scala 31:69:@43262.4]
  assign _T_99973 = portQ_15 ? 16'h400 : _T_99972; // @[Mux.scala 31:69:@43263.4]
  assign _T_99974 = portQ_14 ? 16'h200 : _T_99973; // @[Mux.scala 31:69:@43264.4]
  assign _T_99975 = portQ_13 ? 16'h100 : _T_99974; // @[Mux.scala 31:69:@43265.4]
  assign _T_99976 = portQ_12 ? 16'h80 : _T_99975; // @[Mux.scala 31:69:@43266.4]
  assign _T_99977 = portQ_11 ? 16'h40 : _T_99976; // @[Mux.scala 31:69:@43267.4]
  assign _T_99978 = portQ_10 ? 16'h20 : _T_99977; // @[Mux.scala 31:69:@43268.4]
  assign _T_99979 = portQ_9 ? 16'h10 : _T_99978; // @[Mux.scala 31:69:@43269.4]
  assign _T_99980 = portQ_8 ? 16'h8 : _T_99979; // @[Mux.scala 31:69:@43270.4]
  assign _T_99981 = portQ_7 ? 16'h4 : _T_99980; // @[Mux.scala 31:69:@43271.4]
  assign _T_99982 = portQ_6 ? 16'h2 : _T_99981; // @[Mux.scala 31:69:@43272.4]
  assign _T_99983 = portQ_5 ? 16'h1 : _T_99982; // @[Mux.scala 31:69:@43273.4]
  assign _T_99984 = _T_99983[0]; // @[OneHot.scala 66:30:@43274.4]
  assign _T_99985 = _T_99983[1]; // @[OneHot.scala 66:30:@43275.4]
  assign _T_99986 = _T_99983[2]; // @[OneHot.scala 66:30:@43276.4]
  assign _T_99987 = _T_99983[3]; // @[OneHot.scala 66:30:@43277.4]
  assign _T_99988 = _T_99983[4]; // @[OneHot.scala 66:30:@43278.4]
  assign _T_99989 = _T_99983[5]; // @[OneHot.scala 66:30:@43279.4]
  assign _T_99990 = _T_99983[6]; // @[OneHot.scala 66:30:@43280.4]
  assign _T_99991 = _T_99983[7]; // @[OneHot.scala 66:30:@43281.4]
  assign _T_99992 = _T_99983[8]; // @[OneHot.scala 66:30:@43282.4]
  assign _T_99993 = _T_99983[9]; // @[OneHot.scala 66:30:@43283.4]
  assign _T_99994 = _T_99983[10]; // @[OneHot.scala 66:30:@43284.4]
  assign _T_99995 = _T_99983[11]; // @[OneHot.scala 66:30:@43285.4]
  assign _T_99996 = _T_99983[12]; // @[OneHot.scala 66:30:@43286.4]
  assign _T_99997 = _T_99983[13]; // @[OneHot.scala 66:30:@43287.4]
  assign _T_99998 = _T_99983[14]; // @[OneHot.scala 66:30:@43288.4]
  assign _T_99999 = _T_99983[15]; // @[OneHot.scala 66:30:@43289.4]
  assign _T_100040 = portQ_5 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43307.4]
  assign _T_100041 = portQ_4 ? 16'h4000 : _T_100040; // @[Mux.scala 31:69:@43308.4]
  assign _T_100042 = portQ_3 ? 16'h2000 : _T_100041; // @[Mux.scala 31:69:@43309.4]
  assign _T_100043 = portQ_2 ? 16'h1000 : _T_100042; // @[Mux.scala 31:69:@43310.4]
  assign _T_100044 = portQ_1 ? 16'h800 : _T_100043; // @[Mux.scala 31:69:@43311.4]
  assign _T_100045 = portQ_0 ? 16'h400 : _T_100044; // @[Mux.scala 31:69:@43312.4]
  assign _T_100046 = portQ_15 ? 16'h200 : _T_100045; // @[Mux.scala 31:69:@43313.4]
  assign _T_100047 = portQ_14 ? 16'h100 : _T_100046; // @[Mux.scala 31:69:@43314.4]
  assign _T_100048 = portQ_13 ? 16'h80 : _T_100047; // @[Mux.scala 31:69:@43315.4]
  assign _T_100049 = portQ_12 ? 16'h40 : _T_100048; // @[Mux.scala 31:69:@43316.4]
  assign _T_100050 = portQ_11 ? 16'h20 : _T_100049; // @[Mux.scala 31:69:@43317.4]
  assign _T_100051 = portQ_10 ? 16'h10 : _T_100050; // @[Mux.scala 31:69:@43318.4]
  assign _T_100052 = portQ_9 ? 16'h8 : _T_100051; // @[Mux.scala 31:69:@43319.4]
  assign _T_100053 = portQ_8 ? 16'h4 : _T_100052; // @[Mux.scala 31:69:@43320.4]
  assign _T_100054 = portQ_7 ? 16'h2 : _T_100053; // @[Mux.scala 31:69:@43321.4]
  assign _T_100055 = portQ_6 ? 16'h1 : _T_100054; // @[Mux.scala 31:69:@43322.4]
  assign _T_100056 = _T_100055[0]; // @[OneHot.scala 66:30:@43323.4]
  assign _T_100057 = _T_100055[1]; // @[OneHot.scala 66:30:@43324.4]
  assign _T_100058 = _T_100055[2]; // @[OneHot.scala 66:30:@43325.4]
  assign _T_100059 = _T_100055[3]; // @[OneHot.scala 66:30:@43326.4]
  assign _T_100060 = _T_100055[4]; // @[OneHot.scala 66:30:@43327.4]
  assign _T_100061 = _T_100055[5]; // @[OneHot.scala 66:30:@43328.4]
  assign _T_100062 = _T_100055[6]; // @[OneHot.scala 66:30:@43329.4]
  assign _T_100063 = _T_100055[7]; // @[OneHot.scala 66:30:@43330.4]
  assign _T_100064 = _T_100055[8]; // @[OneHot.scala 66:30:@43331.4]
  assign _T_100065 = _T_100055[9]; // @[OneHot.scala 66:30:@43332.4]
  assign _T_100066 = _T_100055[10]; // @[OneHot.scala 66:30:@43333.4]
  assign _T_100067 = _T_100055[11]; // @[OneHot.scala 66:30:@43334.4]
  assign _T_100068 = _T_100055[12]; // @[OneHot.scala 66:30:@43335.4]
  assign _T_100069 = _T_100055[13]; // @[OneHot.scala 66:30:@43336.4]
  assign _T_100070 = _T_100055[14]; // @[OneHot.scala 66:30:@43337.4]
  assign _T_100071 = _T_100055[15]; // @[OneHot.scala 66:30:@43338.4]
  assign _T_100112 = portQ_6 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43356.4]
  assign _T_100113 = portQ_5 ? 16'h4000 : _T_100112; // @[Mux.scala 31:69:@43357.4]
  assign _T_100114 = portQ_4 ? 16'h2000 : _T_100113; // @[Mux.scala 31:69:@43358.4]
  assign _T_100115 = portQ_3 ? 16'h1000 : _T_100114; // @[Mux.scala 31:69:@43359.4]
  assign _T_100116 = portQ_2 ? 16'h800 : _T_100115; // @[Mux.scala 31:69:@43360.4]
  assign _T_100117 = portQ_1 ? 16'h400 : _T_100116; // @[Mux.scala 31:69:@43361.4]
  assign _T_100118 = portQ_0 ? 16'h200 : _T_100117; // @[Mux.scala 31:69:@43362.4]
  assign _T_100119 = portQ_15 ? 16'h100 : _T_100118; // @[Mux.scala 31:69:@43363.4]
  assign _T_100120 = portQ_14 ? 16'h80 : _T_100119; // @[Mux.scala 31:69:@43364.4]
  assign _T_100121 = portQ_13 ? 16'h40 : _T_100120; // @[Mux.scala 31:69:@43365.4]
  assign _T_100122 = portQ_12 ? 16'h20 : _T_100121; // @[Mux.scala 31:69:@43366.4]
  assign _T_100123 = portQ_11 ? 16'h10 : _T_100122; // @[Mux.scala 31:69:@43367.4]
  assign _T_100124 = portQ_10 ? 16'h8 : _T_100123; // @[Mux.scala 31:69:@43368.4]
  assign _T_100125 = portQ_9 ? 16'h4 : _T_100124; // @[Mux.scala 31:69:@43369.4]
  assign _T_100126 = portQ_8 ? 16'h2 : _T_100125; // @[Mux.scala 31:69:@43370.4]
  assign _T_100127 = portQ_7 ? 16'h1 : _T_100126; // @[Mux.scala 31:69:@43371.4]
  assign _T_100128 = _T_100127[0]; // @[OneHot.scala 66:30:@43372.4]
  assign _T_100129 = _T_100127[1]; // @[OneHot.scala 66:30:@43373.4]
  assign _T_100130 = _T_100127[2]; // @[OneHot.scala 66:30:@43374.4]
  assign _T_100131 = _T_100127[3]; // @[OneHot.scala 66:30:@43375.4]
  assign _T_100132 = _T_100127[4]; // @[OneHot.scala 66:30:@43376.4]
  assign _T_100133 = _T_100127[5]; // @[OneHot.scala 66:30:@43377.4]
  assign _T_100134 = _T_100127[6]; // @[OneHot.scala 66:30:@43378.4]
  assign _T_100135 = _T_100127[7]; // @[OneHot.scala 66:30:@43379.4]
  assign _T_100136 = _T_100127[8]; // @[OneHot.scala 66:30:@43380.4]
  assign _T_100137 = _T_100127[9]; // @[OneHot.scala 66:30:@43381.4]
  assign _T_100138 = _T_100127[10]; // @[OneHot.scala 66:30:@43382.4]
  assign _T_100139 = _T_100127[11]; // @[OneHot.scala 66:30:@43383.4]
  assign _T_100140 = _T_100127[12]; // @[OneHot.scala 66:30:@43384.4]
  assign _T_100141 = _T_100127[13]; // @[OneHot.scala 66:30:@43385.4]
  assign _T_100142 = _T_100127[14]; // @[OneHot.scala 66:30:@43386.4]
  assign _T_100143 = _T_100127[15]; // @[OneHot.scala 66:30:@43387.4]
  assign _T_100184 = portQ_7 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43405.4]
  assign _T_100185 = portQ_6 ? 16'h4000 : _T_100184; // @[Mux.scala 31:69:@43406.4]
  assign _T_100186 = portQ_5 ? 16'h2000 : _T_100185; // @[Mux.scala 31:69:@43407.4]
  assign _T_100187 = portQ_4 ? 16'h1000 : _T_100186; // @[Mux.scala 31:69:@43408.4]
  assign _T_100188 = portQ_3 ? 16'h800 : _T_100187; // @[Mux.scala 31:69:@43409.4]
  assign _T_100189 = portQ_2 ? 16'h400 : _T_100188; // @[Mux.scala 31:69:@43410.4]
  assign _T_100190 = portQ_1 ? 16'h200 : _T_100189; // @[Mux.scala 31:69:@43411.4]
  assign _T_100191 = portQ_0 ? 16'h100 : _T_100190; // @[Mux.scala 31:69:@43412.4]
  assign _T_100192 = portQ_15 ? 16'h80 : _T_100191; // @[Mux.scala 31:69:@43413.4]
  assign _T_100193 = portQ_14 ? 16'h40 : _T_100192; // @[Mux.scala 31:69:@43414.4]
  assign _T_100194 = portQ_13 ? 16'h20 : _T_100193; // @[Mux.scala 31:69:@43415.4]
  assign _T_100195 = portQ_12 ? 16'h10 : _T_100194; // @[Mux.scala 31:69:@43416.4]
  assign _T_100196 = portQ_11 ? 16'h8 : _T_100195; // @[Mux.scala 31:69:@43417.4]
  assign _T_100197 = portQ_10 ? 16'h4 : _T_100196; // @[Mux.scala 31:69:@43418.4]
  assign _T_100198 = portQ_9 ? 16'h2 : _T_100197; // @[Mux.scala 31:69:@43419.4]
  assign _T_100199 = portQ_8 ? 16'h1 : _T_100198; // @[Mux.scala 31:69:@43420.4]
  assign _T_100200 = _T_100199[0]; // @[OneHot.scala 66:30:@43421.4]
  assign _T_100201 = _T_100199[1]; // @[OneHot.scala 66:30:@43422.4]
  assign _T_100202 = _T_100199[2]; // @[OneHot.scala 66:30:@43423.4]
  assign _T_100203 = _T_100199[3]; // @[OneHot.scala 66:30:@43424.4]
  assign _T_100204 = _T_100199[4]; // @[OneHot.scala 66:30:@43425.4]
  assign _T_100205 = _T_100199[5]; // @[OneHot.scala 66:30:@43426.4]
  assign _T_100206 = _T_100199[6]; // @[OneHot.scala 66:30:@43427.4]
  assign _T_100207 = _T_100199[7]; // @[OneHot.scala 66:30:@43428.4]
  assign _T_100208 = _T_100199[8]; // @[OneHot.scala 66:30:@43429.4]
  assign _T_100209 = _T_100199[9]; // @[OneHot.scala 66:30:@43430.4]
  assign _T_100210 = _T_100199[10]; // @[OneHot.scala 66:30:@43431.4]
  assign _T_100211 = _T_100199[11]; // @[OneHot.scala 66:30:@43432.4]
  assign _T_100212 = _T_100199[12]; // @[OneHot.scala 66:30:@43433.4]
  assign _T_100213 = _T_100199[13]; // @[OneHot.scala 66:30:@43434.4]
  assign _T_100214 = _T_100199[14]; // @[OneHot.scala 66:30:@43435.4]
  assign _T_100215 = _T_100199[15]; // @[OneHot.scala 66:30:@43436.4]
  assign _T_100256 = portQ_8 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43454.4]
  assign _T_100257 = portQ_7 ? 16'h4000 : _T_100256; // @[Mux.scala 31:69:@43455.4]
  assign _T_100258 = portQ_6 ? 16'h2000 : _T_100257; // @[Mux.scala 31:69:@43456.4]
  assign _T_100259 = portQ_5 ? 16'h1000 : _T_100258; // @[Mux.scala 31:69:@43457.4]
  assign _T_100260 = portQ_4 ? 16'h800 : _T_100259; // @[Mux.scala 31:69:@43458.4]
  assign _T_100261 = portQ_3 ? 16'h400 : _T_100260; // @[Mux.scala 31:69:@43459.4]
  assign _T_100262 = portQ_2 ? 16'h200 : _T_100261; // @[Mux.scala 31:69:@43460.4]
  assign _T_100263 = portQ_1 ? 16'h100 : _T_100262; // @[Mux.scala 31:69:@43461.4]
  assign _T_100264 = portQ_0 ? 16'h80 : _T_100263; // @[Mux.scala 31:69:@43462.4]
  assign _T_100265 = portQ_15 ? 16'h40 : _T_100264; // @[Mux.scala 31:69:@43463.4]
  assign _T_100266 = portQ_14 ? 16'h20 : _T_100265; // @[Mux.scala 31:69:@43464.4]
  assign _T_100267 = portQ_13 ? 16'h10 : _T_100266; // @[Mux.scala 31:69:@43465.4]
  assign _T_100268 = portQ_12 ? 16'h8 : _T_100267; // @[Mux.scala 31:69:@43466.4]
  assign _T_100269 = portQ_11 ? 16'h4 : _T_100268; // @[Mux.scala 31:69:@43467.4]
  assign _T_100270 = portQ_10 ? 16'h2 : _T_100269; // @[Mux.scala 31:69:@43468.4]
  assign _T_100271 = portQ_9 ? 16'h1 : _T_100270; // @[Mux.scala 31:69:@43469.4]
  assign _T_100272 = _T_100271[0]; // @[OneHot.scala 66:30:@43470.4]
  assign _T_100273 = _T_100271[1]; // @[OneHot.scala 66:30:@43471.4]
  assign _T_100274 = _T_100271[2]; // @[OneHot.scala 66:30:@43472.4]
  assign _T_100275 = _T_100271[3]; // @[OneHot.scala 66:30:@43473.4]
  assign _T_100276 = _T_100271[4]; // @[OneHot.scala 66:30:@43474.4]
  assign _T_100277 = _T_100271[5]; // @[OneHot.scala 66:30:@43475.4]
  assign _T_100278 = _T_100271[6]; // @[OneHot.scala 66:30:@43476.4]
  assign _T_100279 = _T_100271[7]; // @[OneHot.scala 66:30:@43477.4]
  assign _T_100280 = _T_100271[8]; // @[OneHot.scala 66:30:@43478.4]
  assign _T_100281 = _T_100271[9]; // @[OneHot.scala 66:30:@43479.4]
  assign _T_100282 = _T_100271[10]; // @[OneHot.scala 66:30:@43480.4]
  assign _T_100283 = _T_100271[11]; // @[OneHot.scala 66:30:@43481.4]
  assign _T_100284 = _T_100271[12]; // @[OneHot.scala 66:30:@43482.4]
  assign _T_100285 = _T_100271[13]; // @[OneHot.scala 66:30:@43483.4]
  assign _T_100286 = _T_100271[14]; // @[OneHot.scala 66:30:@43484.4]
  assign _T_100287 = _T_100271[15]; // @[OneHot.scala 66:30:@43485.4]
  assign _T_100328 = portQ_9 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43503.4]
  assign _T_100329 = portQ_8 ? 16'h4000 : _T_100328; // @[Mux.scala 31:69:@43504.4]
  assign _T_100330 = portQ_7 ? 16'h2000 : _T_100329; // @[Mux.scala 31:69:@43505.4]
  assign _T_100331 = portQ_6 ? 16'h1000 : _T_100330; // @[Mux.scala 31:69:@43506.4]
  assign _T_100332 = portQ_5 ? 16'h800 : _T_100331; // @[Mux.scala 31:69:@43507.4]
  assign _T_100333 = portQ_4 ? 16'h400 : _T_100332; // @[Mux.scala 31:69:@43508.4]
  assign _T_100334 = portQ_3 ? 16'h200 : _T_100333; // @[Mux.scala 31:69:@43509.4]
  assign _T_100335 = portQ_2 ? 16'h100 : _T_100334; // @[Mux.scala 31:69:@43510.4]
  assign _T_100336 = portQ_1 ? 16'h80 : _T_100335; // @[Mux.scala 31:69:@43511.4]
  assign _T_100337 = portQ_0 ? 16'h40 : _T_100336; // @[Mux.scala 31:69:@43512.4]
  assign _T_100338 = portQ_15 ? 16'h20 : _T_100337; // @[Mux.scala 31:69:@43513.4]
  assign _T_100339 = portQ_14 ? 16'h10 : _T_100338; // @[Mux.scala 31:69:@43514.4]
  assign _T_100340 = portQ_13 ? 16'h8 : _T_100339; // @[Mux.scala 31:69:@43515.4]
  assign _T_100341 = portQ_12 ? 16'h4 : _T_100340; // @[Mux.scala 31:69:@43516.4]
  assign _T_100342 = portQ_11 ? 16'h2 : _T_100341; // @[Mux.scala 31:69:@43517.4]
  assign _T_100343 = portQ_10 ? 16'h1 : _T_100342; // @[Mux.scala 31:69:@43518.4]
  assign _T_100344 = _T_100343[0]; // @[OneHot.scala 66:30:@43519.4]
  assign _T_100345 = _T_100343[1]; // @[OneHot.scala 66:30:@43520.4]
  assign _T_100346 = _T_100343[2]; // @[OneHot.scala 66:30:@43521.4]
  assign _T_100347 = _T_100343[3]; // @[OneHot.scala 66:30:@43522.4]
  assign _T_100348 = _T_100343[4]; // @[OneHot.scala 66:30:@43523.4]
  assign _T_100349 = _T_100343[5]; // @[OneHot.scala 66:30:@43524.4]
  assign _T_100350 = _T_100343[6]; // @[OneHot.scala 66:30:@43525.4]
  assign _T_100351 = _T_100343[7]; // @[OneHot.scala 66:30:@43526.4]
  assign _T_100352 = _T_100343[8]; // @[OneHot.scala 66:30:@43527.4]
  assign _T_100353 = _T_100343[9]; // @[OneHot.scala 66:30:@43528.4]
  assign _T_100354 = _T_100343[10]; // @[OneHot.scala 66:30:@43529.4]
  assign _T_100355 = _T_100343[11]; // @[OneHot.scala 66:30:@43530.4]
  assign _T_100356 = _T_100343[12]; // @[OneHot.scala 66:30:@43531.4]
  assign _T_100357 = _T_100343[13]; // @[OneHot.scala 66:30:@43532.4]
  assign _T_100358 = _T_100343[14]; // @[OneHot.scala 66:30:@43533.4]
  assign _T_100359 = _T_100343[15]; // @[OneHot.scala 66:30:@43534.4]
  assign _T_100400 = portQ_10 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43552.4]
  assign _T_100401 = portQ_9 ? 16'h4000 : _T_100400; // @[Mux.scala 31:69:@43553.4]
  assign _T_100402 = portQ_8 ? 16'h2000 : _T_100401; // @[Mux.scala 31:69:@43554.4]
  assign _T_100403 = portQ_7 ? 16'h1000 : _T_100402; // @[Mux.scala 31:69:@43555.4]
  assign _T_100404 = portQ_6 ? 16'h800 : _T_100403; // @[Mux.scala 31:69:@43556.4]
  assign _T_100405 = portQ_5 ? 16'h400 : _T_100404; // @[Mux.scala 31:69:@43557.4]
  assign _T_100406 = portQ_4 ? 16'h200 : _T_100405; // @[Mux.scala 31:69:@43558.4]
  assign _T_100407 = portQ_3 ? 16'h100 : _T_100406; // @[Mux.scala 31:69:@43559.4]
  assign _T_100408 = portQ_2 ? 16'h80 : _T_100407; // @[Mux.scala 31:69:@43560.4]
  assign _T_100409 = portQ_1 ? 16'h40 : _T_100408; // @[Mux.scala 31:69:@43561.4]
  assign _T_100410 = portQ_0 ? 16'h20 : _T_100409; // @[Mux.scala 31:69:@43562.4]
  assign _T_100411 = portQ_15 ? 16'h10 : _T_100410; // @[Mux.scala 31:69:@43563.4]
  assign _T_100412 = portQ_14 ? 16'h8 : _T_100411; // @[Mux.scala 31:69:@43564.4]
  assign _T_100413 = portQ_13 ? 16'h4 : _T_100412; // @[Mux.scala 31:69:@43565.4]
  assign _T_100414 = portQ_12 ? 16'h2 : _T_100413; // @[Mux.scala 31:69:@43566.4]
  assign _T_100415 = portQ_11 ? 16'h1 : _T_100414; // @[Mux.scala 31:69:@43567.4]
  assign _T_100416 = _T_100415[0]; // @[OneHot.scala 66:30:@43568.4]
  assign _T_100417 = _T_100415[1]; // @[OneHot.scala 66:30:@43569.4]
  assign _T_100418 = _T_100415[2]; // @[OneHot.scala 66:30:@43570.4]
  assign _T_100419 = _T_100415[3]; // @[OneHot.scala 66:30:@43571.4]
  assign _T_100420 = _T_100415[4]; // @[OneHot.scala 66:30:@43572.4]
  assign _T_100421 = _T_100415[5]; // @[OneHot.scala 66:30:@43573.4]
  assign _T_100422 = _T_100415[6]; // @[OneHot.scala 66:30:@43574.4]
  assign _T_100423 = _T_100415[7]; // @[OneHot.scala 66:30:@43575.4]
  assign _T_100424 = _T_100415[8]; // @[OneHot.scala 66:30:@43576.4]
  assign _T_100425 = _T_100415[9]; // @[OneHot.scala 66:30:@43577.4]
  assign _T_100426 = _T_100415[10]; // @[OneHot.scala 66:30:@43578.4]
  assign _T_100427 = _T_100415[11]; // @[OneHot.scala 66:30:@43579.4]
  assign _T_100428 = _T_100415[12]; // @[OneHot.scala 66:30:@43580.4]
  assign _T_100429 = _T_100415[13]; // @[OneHot.scala 66:30:@43581.4]
  assign _T_100430 = _T_100415[14]; // @[OneHot.scala 66:30:@43582.4]
  assign _T_100431 = _T_100415[15]; // @[OneHot.scala 66:30:@43583.4]
  assign _T_100472 = portQ_11 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43601.4]
  assign _T_100473 = portQ_10 ? 16'h4000 : _T_100472; // @[Mux.scala 31:69:@43602.4]
  assign _T_100474 = portQ_9 ? 16'h2000 : _T_100473; // @[Mux.scala 31:69:@43603.4]
  assign _T_100475 = portQ_8 ? 16'h1000 : _T_100474; // @[Mux.scala 31:69:@43604.4]
  assign _T_100476 = portQ_7 ? 16'h800 : _T_100475; // @[Mux.scala 31:69:@43605.4]
  assign _T_100477 = portQ_6 ? 16'h400 : _T_100476; // @[Mux.scala 31:69:@43606.4]
  assign _T_100478 = portQ_5 ? 16'h200 : _T_100477; // @[Mux.scala 31:69:@43607.4]
  assign _T_100479 = portQ_4 ? 16'h100 : _T_100478; // @[Mux.scala 31:69:@43608.4]
  assign _T_100480 = portQ_3 ? 16'h80 : _T_100479; // @[Mux.scala 31:69:@43609.4]
  assign _T_100481 = portQ_2 ? 16'h40 : _T_100480; // @[Mux.scala 31:69:@43610.4]
  assign _T_100482 = portQ_1 ? 16'h20 : _T_100481; // @[Mux.scala 31:69:@43611.4]
  assign _T_100483 = portQ_0 ? 16'h10 : _T_100482; // @[Mux.scala 31:69:@43612.4]
  assign _T_100484 = portQ_15 ? 16'h8 : _T_100483; // @[Mux.scala 31:69:@43613.4]
  assign _T_100485 = portQ_14 ? 16'h4 : _T_100484; // @[Mux.scala 31:69:@43614.4]
  assign _T_100486 = portQ_13 ? 16'h2 : _T_100485; // @[Mux.scala 31:69:@43615.4]
  assign _T_100487 = portQ_12 ? 16'h1 : _T_100486; // @[Mux.scala 31:69:@43616.4]
  assign _T_100488 = _T_100487[0]; // @[OneHot.scala 66:30:@43617.4]
  assign _T_100489 = _T_100487[1]; // @[OneHot.scala 66:30:@43618.4]
  assign _T_100490 = _T_100487[2]; // @[OneHot.scala 66:30:@43619.4]
  assign _T_100491 = _T_100487[3]; // @[OneHot.scala 66:30:@43620.4]
  assign _T_100492 = _T_100487[4]; // @[OneHot.scala 66:30:@43621.4]
  assign _T_100493 = _T_100487[5]; // @[OneHot.scala 66:30:@43622.4]
  assign _T_100494 = _T_100487[6]; // @[OneHot.scala 66:30:@43623.4]
  assign _T_100495 = _T_100487[7]; // @[OneHot.scala 66:30:@43624.4]
  assign _T_100496 = _T_100487[8]; // @[OneHot.scala 66:30:@43625.4]
  assign _T_100497 = _T_100487[9]; // @[OneHot.scala 66:30:@43626.4]
  assign _T_100498 = _T_100487[10]; // @[OneHot.scala 66:30:@43627.4]
  assign _T_100499 = _T_100487[11]; // @[OneHot.scala 66:30:@43628.4]
  assign _T_100500 = _T_100487[12]; // @[OneHot.scala 66:30:@43629.4]
  assign _T_100501 = _T_100487[13]; // @[OneHot.scala 66:30:@43630.4]
  assign _T_100502 = _T_100487[14]; // @[OneHot.scala 66:30:@43631.4]
  assign _T_100503 = _T_100487[15]; // @[OneHot.scala 66:30:@43632.4]
  assign _T_100544 = portQ_12 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43650.4]
  assign _T_100545 = portQ_11 ? 16'h4000 : _T_100544; // @[Mux.scala 31:69:@43651.4]
  assign _T_100546 = portQ_10 ? 16'h2000 : _T_100545; // @[Mux.scala 31:69:@43652.4]
  assign _T_100547 = portQ_9 ? 16'h1000 : _T_100546; // @[Mux.scala 31:69:@43653.4]
  assign _T_100548 = portQ_8 ? 16'h800 : _T_100547; // @[Mux.scala 31:69:@43654.4]
  assign _T_100549 = portQ_7 ? 16'h400 : _T_100548; // @[Mux.scala 31:69:@43655.4]
  assign _T_100550 = portQ_6 ? 16'h200 : _T_100549; // @[Mux.scala 31:69:@43656.4]
  assign _T_100551 = portQ_5 ? 16'h100 : _T_100550; // @[Mux.scala 31:69:@43657.4]
  assign _T_100552 = portQ_4 ? 16'h80 : _T_100551; // @[Mux.scala 31:69:@43658.4]
  assign _T_100553 = portQ_3 ? 16'h40 : _T_100552; // @[Mux.scala 31:69:@43659.4]
  assign _T_100554 = portQ_2 ? 16'h20 : _T_100553; // @[Mux.scala 31:69:@43660.4]
  assign _T_100555 = portQ_1 ? 16'h10 : _T_100554; // @[Mux.scala 31:69:@43661.4]
  assign _T_100556 = portQ_0 ? 16'h8 : _T_100555; // @[Mux.scala 31:69:@43662.4]
  assign _T_100557 = portQ_15 ? 16'h4 : _T_100556; // @[Mux.scala 31:69:@43663.4]
  assign _T_100558 = portQ_14 ? 16'h2 : _T_100557; // @[Mux.scala 31:69:@43664.4]
  assign _T_100559 = portQ_13 ? 16'h1 : _T_100558; // @[Mux.scala 31:69:@43665.4]
  assign _T_100560 = _T_100559[0]; // @[OneHot.scala 66:30:@43666.4]
  assign _T_100561 = _T_100559[1]; // @[OneHot.scala 66:30:@43667.4]
  assign _T_100562 = _T_100559[2]; // @[OneHot.scala 66:30:@43668.4]
  assign _T_100563 = _T_100559[3]; // @[OneHot.scala 66:30:@43669.4]
  assign _T_100564 = _T_100559[4]; // @[OneHot.scala 66:30:@43670.4]
  assign _T_100565 = _T_100559[5]; // @[OneHot.scala 66:30:@43671.4]
  assign _T_100566 = _T_100559[6]; // @[OneHot.scala 66:30:@43672.4]
  assign _T_100567 = _T_100559[7]; // @[OneHot.scala 66:30:@43673.4]
  assign _T_100568 = _T_100559[8]; // @[OneHot.scala 66:30:@43674.4]
  assign _T_100569 = _T_100559[9]; // @[OneHot.scala 66:30:@43675.4]
  assign _T_100570 = _T_100559[10]; // @[OneHot.scala 66:30:@43676.4]
  assign _T_100571 = _T_100559[11]; // @[OneHot.scala 66:30:@43677.4]
  assign _T_100572 = _T_100559[12]; // @[OneHot.scala 66:30:@43678.4]
  assign _T_100573 = _T_100559[13]; // @[OneHot.scala 66:30:@43679.4]
  assign _T_100574 = _T_100559[14]; // @[OneHot.scala 66:30:@43680.4]
  assign _T_100575 = _T_100559[15]; // @[OneHot.scala 66:30:@43681.4]
  assign _T_100616 = portQ_13 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43699.4]
  assign _T_100617 = portQ_12 ? 16'h4000 : _T_100616; // @[Mux.scala 31:69:@43700.4]
  assign _T_100618 = portQ_11 ? 16'h2000 : _T_100617; // @[Mux.scala 31:69:@43701.4]
  assign _T_100619 = portQ_10 ? 16'h1000 : _T_100618; // @[Mux.scala 31:69:@43702.4]
  assign _T_100620 = portQ_9 ? 16'h800 : _T_100619; // @[Mux.scala 31:69:@43703.4]
  assign _T_100621 = portQ_8 ? 16'h400 : _T_100620; // @[Mux.scala 31:69:@43704.4]
  assign _T_100622 = portQ_7 ? 16'h200 : _T_100621; // @[Mux.scala 31:69:@43705.4]
  assign _T_100623 = portQ_6 ? 16'h100 : _T_100622; // @[Mux.scala 31:69:@43706.4]
  assign _T_100624 = portQ_5 ? 16'h80 : _T_100623; // @[Mux.scala 31:69:@43707.4]
  assign _T_100625 = portQ_4 ? 16'h40 : _T_100624; // @[Mux.scala 31:69:@43708.4]
  assign _T_100626 = portQ_3 ? 16'h20 : _T_100625; // @[Mux.scala 31:69:@43709.4]
  assign _T_100627 = portQ_2 ? 16'h10 : _T_100626; // @[Mux.scala 31:69:@43710.4]
  assign _T_100628 = portQ_1 ? 16'h8 : _T_100627; // @[Mux.scala 31:69:@43711.4]
  assign _T_100629 = portQ_0 ? 16'h4 : _T_100628; // @[Mux.scala 31:69:@43712.4]
  assign _T_100630 = portQ_15 ? 16'h2 : _T_100629; // @[Mux.scala 31:69:@43713.4]
  assign _T_100631 = portQ_14 ? 16'h1 : _T_100630; // @[Mux.scala 31:69:@43714.4]
  assign _T_100632 = _T_100631[0]; // @[OneHot.scala 66:30:@43715.4]
  assign _T_100633 = _T_100631[1]; // @[OneHot.scala 66:30:@43716.4]
  assign _T_100634 = _T_100631[2]; // @[OneHot.scala 66:30:@43717.4]
  assign _T_100635 = _T_100631[3]; // @[OneHot.scala 66:30:@43718.4]
  assign _T_100636 = _T_100631[4]; // @[OneHot.scala 66:30:@43719.4]
  assign _T_100637 = _T_100631[5]; // @[OneHot.scala 66:30:@43720.4]
  assign _T_100638 = _T_100631[6]; // @[OneHot.scala 66:30:@43721.4]
  assign _T_100639 = _T_100631[7]; // @[OneHot.scala 66:30:@43722.4]
  assign _T_100640 = _T_100631[8]; // @[OneHot.scala 66:30:@43723.4]
  assign _T_100641 = _T_100631[9]; // @[OneHot.scala 66:30:@43724.4]
  assign _T_100642 = _T_100631[10]; // @[OneHot.scala 66:30:@43725.4]
  assign _T_100643 = _T_100631[11]; // @[OneHot.scala 66:30:@43726.4]
  assign _T_100644 = _T_100631[12]; // @[OneHot.scala 66:30:@43727.4]
  assign _T_100645 = _T_100631[13]; // @[OneHot.scala 66:30:@43728.4]
  assign _T_100646 = _T_100631[14]; // @[OneHot.scala 66:30:@43729.4]
  assign _T_100647 = _T_100631[15]; // @[OneHot.scala 66:30:@43730.4]
  assign _T_100688 = portQ_14 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43748.4]
  assign _T_100689 = portQ_13 ? 16'h4000 : _T_100688; // @[Mux.scala 31:69:@43749.4]
  assign _T_100690 = portQ_12 ? 16'h2000 : _T_100689; // @[Mux.scala 31:69:@43750.4]
  assign _T_100691 = portQ_11 ? 16'h1000 : _T_100690; // @[Mux.scala 31:69:@43751.4]
  assign _T_100692 = portQ_10 ? 16'h800 : _T_100691; // @[Mux.scala 31:69:@43752.4]
  assign _T_100693 = portQ_9 ? 16'h400 : _T_100692; // @[Mux.scala 31:69:@43753.4]
  assign _T_100694 = portQ_8 ? 16'h200 : _T_100693; // @[Mux.scala 31:69:@43754.4]
  assign _T_100695 = portQ_7 ? 16'h100 : _T_100694; // @[Mux.scala 31:69:@43755.4]
  assign _T_100696 = portQ_6 ? 16'h80 : _T_100695; // @[Mux.scala 31:69:@43756.4]
  assign _T_100697 = portQ_5 ? 16'h40 : _T_100696; // @[Mux.scala 31:69:@43757.4]
  assign _T_100698 = portQ_4 ? 16'h20 : _T_100697; // @[Mux.scala 31:69:@43758.4]
  assign _T_100699 = portQ_3 ? 16'h10 : _T_100698; // @[Mux.scala 31:69:@43759.4]
  assign _T_100700 = portQ_2 ? 16'h8 : _T_100699; // @[Mux.scala 31:69:@43760.4]
  assign _T_100701 = portQ_1 ? 16'h4 : _T_100700; // @[Mux.scala 31:69:@43761.4]
  assign _T_100702 = portQ_0 ? 16'h2 : _T_100701; // @[Mux.scala 31:69:@43762.4]
  assign _T_100703 = portQ_15 ? 16'h1 : _T_100702; // @[Mux.scala 31:69:@43763.4]
  assign _T_100704 = _T_100703[0]; // @[OneHot.scala 66:30:@43764.4]
  assign _T_100705 = _T_100703[1]; // @[OneHot.scala 66:30:@43765.4]
  assign _T_100706 = _T_100703[2]; // @[OneHot.scala 66:30:@43766.4]
  assign _T_100707 = _T_100703[3]; // @[OneHot.scala 66:30:@43767.4]
  assign _T_100708 = _T_100703[4]; // @[OneHot.scala 66:30:@43768.4]
  assign _T_100709 = _T_100703[5]; // @[OneHot.scala 66:30:@43769.4]
  assign _T_100710 = _T_100703[6]; // @[OneHot.scala 66:30:@43770.4]
  assign _T_100711 = _T_100703[7]; // @[OneHot.scala 66:30:@43771.4]
  assign _T_100712 = _T_100703[8]; // @[OneHot.scala 66:30:@43772.4]
  assign _T_100713 = _T_100703[9]; // @[OneHot.scala 66:30:@43773.4]
  assign _T_100714 = _T_100703[10]; // @[OneHot.scala 66:30:@43774.4]
  assign _T_100715 = _T_100703[11]; // @[OneHot.scala 66:30:@43775.4]
  assign _T_100716 = _T_100703[12]; // @[OneHot.scala 66:30:@43776.4]
  assign _T_100717 = _T_100703[13]; // @[OneHot.scala 66:30:@43777.4]
  assign _T_100718 = _T_100703[14]; // @[OneHot.scala 66:30:@43778.4]
  assign _T_100719 = _T_100703[15]; // @[OneHot.scala 66:30:@43779.4]
  assign _T_100784 = {_T_99631,_T_99630,_T_99629,_T_99628,_T_99627,_T_99626,_T_99625,_T_99624}; // @[Mux.scala 19:72:@43803.4]
  assign _T_100792 = {_T_99639,_T_99638,_T_99637,_T_99636,_T_99635,_T_99634,_T_99633,_T_99632,_T_100784}; // @[Mux.scala 19:72:@43811.4]
  assign _T_100794 = _T_90408 ? _T_100792 : 16'h0; // @[Mux.scala 19:72:@43812.4]
  assign _T_100801 = {_T_99702,_T_99701,_T_99700,_T_99699,_T_99698,_T_99697,_T_99696,_T_99711}; // @[Mux.scala 19:72:@43819.4]
  assign _T_100809 = {_T_99710,_T_99709,_T_99708,_T_99707,_T_99706,_T_99705,_T_99704,_T_99703,_T_100801}; // @[Mux.scala 19:72:@43827.4]
  assign _T_100811 = _T_90409 ? _T_100809 : 16'h0; // @[Mux.scala 19:72:@43828.4]
  assign _T_100818 = {_T_99773,_T_99772,_T_99771,_T_99770,_T_99769,_T_99768,_T_99783,_T_99782}; // @[Mux.scala 19:72:@43835.4]
  assign _T_100826 = {_T_99781,_T_99780,_T_99779,_T_99778,_T_99777,_T_99776,_T_99775,_T_99774,_T_100818}; // @[Mux.scala 19:72:@43843.4]
  assign _T_100828 = _T_90410 ? _T_100826 : 16'h0; // @[Mux.scala 19:72:@43844.4]
  assign _T_100835 = {_T_99844,_T_99843,_T_99842,_T_99841,_T_99840,_T_99855,_T_99854,_T_99853}; // @[Mux.scala 19:72:@43851.4]
  assign _T_100843 = {_T_99852,_T_99851,_T_99850,_T_99849,_T_99848,_T_99847,_T_99846,_T_99845,_T_100835}; // @[Mux.scala 19:72:@43859.4]
  assign _T_100845 = _T_90411 ? _T_100843 : 16'h0; // @[Mux.scala 19:72:@43860.4]
  assign _T_100852 = {_T_99915,_T_99914,_T_99913,_T_99912,_T_99927,_T_99926,_T_99925,_T_99924}; // @[Mux.scala 19:72:@43867.4]
  assign _T_100860 = {_T_99923,_T_99922,_T_99921,_T_99920,_T_99919,_T_99918,_T_99917,_T_99916,_T_100852}; // @[Mux.scala 19:72:@43875.4]
  assign _T_100862 = _T_90412 ? _T_100860 : 16'h0; // @[Mux.scala 19:72:@43876.4]
  assign _T_100869 = {_T_99986,_T_99985,_T_99984,_T_99999,_T_99998,_T_99997,_T_99996,_T_99995}; // @[Mux.scala 19:72:@43883.4]
  assign _T_100877 = {_T_99994,_T_99993,_T_99992,_T_99991,_T_99990,_T_99989,_T_99988,_T_99987,_T_100869}; // @[Mux.scala 19:72:@43891.4]
  assign _T_100879 = _T_90413 ? _T_100877 : 16'h0; // @[Mux.scala 19:72:@43892.4]
  assign _T_100886 = {_T_100057,_T_100056,_T_100071,_T_100070,_T_100069,_T_100068,_T_100067,_T_100066}; // @[Mux.scala 19:72:@43899.4]
  assign _T_100894 = {_T_100065,_T_100064,_T_100063,_T_100062,_T_100061,_T_100060,_T_100059,_T_100058,_T_100886}; // @[Mux.scala 19:72:@43907.4]
  assign _T_100896 = _T_90414 ? _T_100894 : 16'h0; // @[Mux.scala 19:72:@43908.4]
  assign _T_100903 = {_T_100128,_T_100143,_T_100142,_T_100141,_T_100140,_T_100139,_T_100138,_T_100137}; // @[Mux.scala 19:72:@43915.4]
  assign _T_100911 = {_T_100136,_T_100135,_T_100134,_T_100133,_T_100132,_T_100131,_T_100130,_T_100129,_T_100903}; // @[Mux.scala 19:72:@43923.4]
  assign _T_100913 = _T_90415 ? _T_100911 : 16'h0; // @[Mux.scala 19:72:@43924.4]
  assign _T_100920 = {_T_100215,_T_100214,_T_100213,_T_100212,_T_100211,_T_100210,_T_100209,_T_100208}; // @[Mux.scala 19:72:@43931.4]
  assign _T_100928 = {_T_100207,_T_100206,_T_100205,_T_100204,_T_100203,_T_100202,_T_100201,_T_100200,_T_100920}; // @[Mux.scala 19:72:@43939.4]
  assign _T_100930 = _T_90416 ? _T_100928 : 16'h0; // @[Mux.scala 19:72:@43940.4]
  assign _T_100937 = {_T_100286,_T_100285,_T_100284,_T_100283,_T_100282,_T_100281,_T_100280,_T_100279}; // @[Mux.scala 19:72:@43947.4]
  assign _T_100945 = {_T_100278,_T_100277,_T_100276,_T_100275,_T_100274,_T_100273,_T_100272,_T_100287,_T_100937}; // @[Mux.scala 19:72:@43955.4]
  assign _T_100947 = _T_90417 ? _T_100945 : 16'h0; // @[Mux.scala 19:72:@43956.4]
  assign _T_100954 = {_T_100357,_T_100356,_T_100355,_T_100354,_T_100353,_T_100352,_T_100351,_T_100350}; // @[Mux.scala 19:72:@43963.4]
  assign _T_100962 = {_T_100349,_T_100348,_T_100347,_T_100346,_T_100345,_T_100344,_T_100359,_T_100358,_T_100954}; // @[Mux.scala 19:72:@43971.4]
  assign _T_100964 = _T_90418 ? _T_100962 : 16'h0; // @[Mux.scala 19:72:@43972.4]
  assign _T_100971 = {_T_100428,_T_100427,_T_100426,_T_100425,_T_100424,_T_100423,_T_100422,_T_100421}; // @[Mux.scala 19:72:@43979.4]
  assign _T_100979 = {_T_100420,_T_100419,_T_100418,_T_100417,_T_100416,_T_100431,_T_100430,_T_100429,_T_100971}; // @[Mux.scala 19:72:@43987.4]
  assign _T_100981 = _T_90419 ? _T_100979 : 16'h0; // @[Mux.scala 19:72:@43988.4]
  assign _T_100988 = {_T_100499,_T_100498,_T_100497,_T_100496,_T_100495,_T_100494,_T_100493,_T_100492}; // @[Mux.scala 19:72:@43995.4]
  assign _T_100996 = {_T_100491,_T_100490,_T_100489,_T_100488,_T_100503,_T_100502,_T_100501,_T_100500,_T_100988}; // @[Mux.scala 19:72:@44003.4]
  assign _T_100998 = _T_90420 ? _T_100996 : 16'h0; // @[Mux.scala 19:72:@44004.4]
  assign _T_101005 = {_T_100570,_T_100569,_T_100568,_T_100567,_T_100566,_T_100565,_T_100564,_T_100563}; // @[Mux.scala 19:72:@44011.4]
  assign _T_101013 = {_T_100562,_T_100561,_T_100560,_T_100575,_T_100574,_T_100573,_T_100572,_T_100571,_T_101005}; // @[Mux.scala 19:72:@44019.4]
  assign _T_101015 = _T_90421 ? _T_101013 : 16'h0; // @[Mux.scala 19:72:@44020.4]
  assign _T_101022 = {_T_100641,_T_100640,_T_100639,_T_100638,_T_100637,_T_100636,_T_100635,_T_100634}; // @[Mux.scala 19:72:@44027.4]
  assign _T_101030 = {_T_100633,_T_100632,_T_100647,_T_100646,_T_100645,_T_100644,_T_100643,_T_100642,_T_101022}; // @[Mux.scala 19:72:@44035.4]
  assign _T_101032 = _T_90422 ? _T_101030 : 16'h0; // @[Mux.scala 19:72:@44036.4]
  assign _T_101039 = {_T_100712,_T_100711,_T_100710,_T_100709,_T_100708,_T_100707,_T_100706,_T_100705}; // @[Mux.scala 19:72:@44043.4]
  assign _T_101047 = {_T_100704,_T_100719,_T_100718,_T_100717,_T_100716,_T_100715,_T_100714,_T_100713,_T_101039}; // @[Mux.scala 19:72:@44051.4]
  assign _T_101049 = _T_90423 ? _T_101047 : 16'h0; // @[Mux.scala 19:72:@44052.4]
  assign _T_101050 = _T_100794 | _T_100811; // @[Mux.scala 19:72:@44053.4]
  assign _T_101051 = _T_101050 | _T_100828; // @[Mux.scala 19:72:@44054.4]
  assign _T_101052 = _T_101051 | _T_100845; // @[Mux.scala 19:72:@44055.4]
  assign _T_101053 = _T_101052 | _T_100862; // @[Mux.scala 19:72:@44056.4]
  assign _T_101054 = _T_101053 | _T_100879; // @[Mux.scala 19:72:@44057.4]
  assign _T_101055 = _T_101054 | _T_100896; // @[Mux.scala 19:72:@44058.4]
  assign _T_101056 = _T_101055 | _T_100913; // @[Mux.scala 19:72:@44059.4]
  assign _T_101057 = _T_101056 | _T_100930; // @[Mux.scala 19:72:@44060.4]
  assign _T_101058 = _T_101057 | _T_100947; // @[Mux.scala 19:72:@44061.4]
  assign _T_101059 = _T_101058 | _T_100964; // @[Mux.scala 19:72:@44062.4]
  assign _T_101060 = _T_101059 | _T_100981; // @[Mux.scala 19:72:@44063.4]
  assign _T_101061 = _T_101060 | _T_100998; // @[Mux.scala 19:72:@44064.4]
  assign _T_101062 = _T_101061 | _T_101015; // @[Mux.scala 19:72:@44065.4]
  assign _T_101063 = _T_101062 | _T_101032; // @[Mux.scala 19:72:@44066.4]
  assign _T_101064 = _T_101063 | _T_101049; // @[Mux.scala 19:72:@44067.4]
  assign outputPriorityPorts_1_0 = _T_101064[0]; // @[Mux.scala 19:72:@44071.4]
  assign outputPriorityPorts_1_1 = _T_101064[1]; // @[Mux.scala 19:72:@44073.4]
  assign outputPriorityPorts_1_2 = _T_101064[2]; // @[Mux.scala 19:72:@44075.4]
  assign outputPriorityPorts_1_3 = _T_101064[3]; // @[Mux.scala 19:72:@44077.4]
  assign outputPriorityPorts_1_4 = _T_101064[4]; // @[Mux.scala 19:72:@44079.4]
  assign outputPriorityPorts_1_5 = _T_101064[5]; // @[Mux.scala 19:72:@44081.4]
  assign outputPriorityPorts_1_6 = _T_101064[6]; // @[Mux.scala 19:72:@44083.4]
  assign outputPriorityPorts_1_7 = _T_101064[7]; // @[Mux.scala 19:72:@44085.4]
  assign outputPriorityPorts_1_8 = _T_101064[8]; // @[Mux.scala 19:72:@44087.4]
  assign outputPriorityPorts_1_9 = _T_101064[9]; // @[Mux.scala 19:72:@44089.4]
  assign outputPriorityPorts_1_10 = _T_101064[10]; // @[Mux.scala 19:72:@44091.4]
  assign outputPriorityPorts_1_11 = _T_101064[11]; // @[Mux.scala 19:72:@44093.4]
  assign outputPriorityPorts_1_12 = _T_101064[12]; // @[Mux.scala 19:72:@44095.4]
  assign outputPriorityPorts_1_13 = _T_101064[13]; // @[Mux.scala 19:72:@44097.4]
  assign outputPriorityPorts_1_14 = _T_101064[14]; // @[Mux.scala 19:72:@44099.4]
  assign outputPriorityPorts_1_15 = _T_101064[15]; // @[Mux.scala 19:72:@44101.4]
  assign _T_101207 = inputPriorityPorts_0_0 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44123.6]
  assign _T_101208 = inputPriorityPorts_1_0 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@44124.6]
  assign _T_101219 = _T_101207 | _T_101208; // @[LoadQueue.scala 314:26:@44129.6]
  assign _T_101220 = {_T_101208,_T_101207}; // @[OneHot.scala 18:45:@44131.8]
  assign _T_101221 = _T_101220[1]; // @[CircuitMath.scala 30:8:@44132.8]
  assign _GEN_2115 = _T_101221 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@44133.8]
  assign _GEN_2116 = _T_101219 ? _GEN_2115 : addrQ_0; // @[LoadQueue.scala 314:36:@44130.6]
  assign _GEN_2117 = _T_101219 ? 1'h1 : addrKnown_0; // @[LoadQueue.scala 314:36:@44130.6]
  assign _GEN_2118 = initBits_0 ? 1'h0 : _GEN_2117; // @[LoadQueue.scala 308:34:@44119.4]
  assign _GEN_2119 = initBits_0 ? addrQ_0 : _GEN_2116; // @[LoadQueue.scala 308:34:@44119.4]
  assign _T_101225 = inputPriorityPorts_0_1 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44141.6]
  assign _T_101226 = inputPriorityPorts_1_1 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@44142.6]
  assign _T_101237 = _T_101225 | _T_101226; // @[LoadQueue.scala 314:26:@44147.6]
  assign _T_101238 = {_T_101226,_T_101225}; // @[OneHot.scala 18:45:@44149.8]
  assign _T_101239 = _T_101238[1]; // @[CircuitMath.scala 30:8:@44150.8]
  assign _GEN_2121 = _T_101239 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@44151.8]
  assign _GEN_2122 = _T_101237 ? _GEN_2121 : addrQ_1; // @[LoadQueue.scala 314:36:@44148.6]
  assign _GEN_2123 = _T_101237 ? 1'h1 : addrKnown_1; // @[LoadQueue.scala 314:36:@44148.6]
  assign _GEN_2124 = initBits_1 ? 1'h0 : _GEN_2123; // @[LoadQueue.scala 308:34:@44137.4]
  assign _GEN_2125 = initBits_1 ? addrQ_1 : _GEN_2122; // @[LoadQueue.scala 308:34:@44137.4]
  assign _T_101243 = inputPriorityPorts_0_2 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44159.6]
  assign _T_101244 = inputPriorityPorts_1_2 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@44160.6]
  assign _T_101255 = _T_101243 | _T_101244; // @[LoadQueue.scala 314:26:@44165.6]
  assign _T_101256 = {_T_101244,_T_101243}; // @[OneHot.scala 18:45:@44167.8]
  assign _T_101257 = _T_101256[1]; // @[CircuitMath.scala 30:8:@44168.8]
  assign _GEN_2127 = _T_101257 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@44169.8]
  assign _GEN_2128 = _T_101255 ? _GEN_2127 : addrQ_2; // @[LoadQueue.scala 314:36:@44166.6]
  assign _GEN_2129 = _T_101255 ? 1'h1 : addrKnown_2; // @[LoadQueue.scala 314:36:@44166.6]
  assign _GEN_2130 = initBits_2 ? 1'h0 : _GEN_2129; // @[LoadQueue.scala 308:34:@44155.4]
  assign _GEN_2131 = initBits_2 ? addrQ_2 : _GEN_2128; // @[LoadQueue.scala 308:34:@44155.4]
  assign _T_101261 = inputPriorityPorts_0_3 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44177.6]
  assign _T_101262 = inputPriorityPorts_1_3 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@44178.6]
  assign _T_101273 = _T_101261 | _T_101262; // @[LoadQueue.scala 314:26:@44183.6]
  assign _T_101274 = {_T_101262,_T_101261}; // @[OneHot.scala 18:45:@44185.8]
  assign _T_101275 = _T_101274[1]; // @[CircuitMath.scala 30:8:@44186.8]
  assign _GEN_2133 = _T_101275 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@44187.8]
  assign _GEN_2134 = _T_101273 ? _GEN_2133 : addrQ_3; // @[LoadQueue.scala 314:36:@44184.6]
  assign _GEN_2135 = _T_101273 ? 1'h1 : addrKnown_3; // @[LoadQueue.scala 314:36:@44184.6]
  assign _GEN_2136 = initBits_3 ? 1'h0 : _GEN_2135; // @[LoadQueue.scala 308:34:@44173.4]
  assign _GEN_2137 = initBits_3 ? addrQ_3 : _GEN_2134; // @[LoadQueue.scala 308:34:@44173.4]
  assign _T_101279 = inputPriorityPorts_0_4 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44195.6]
  assign _T_101280 = inputPriorityPorts_1_4 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@44196.6]
  assign _T_101291 = _T_101279 | _T_101280; // @[LoadQueue.scala 314:26:@44201.6]
  assign _T_101292 = {_T_101280,_T_101279}; // @[OneHot.scala 18:45:@44203.8]
  assign _T_101293 = _T_101292[1]; // @[CircuitMath.scala 30:8:@44204.8]
  assign _GEN_2139 = _T_101293 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@44205.8]
  assign _GEN_2140 = _T_101291 ? _GEN_2139 : addrQ_4; // @[LoadQueue.scala 314:36:@44202.6]
  assign _GEN_2141 = _T_101291 ? 1'h1 : addrKnown_4; // @[LoadQueue.scala 314:36:@44202.6]
  assign _GEN_2142 = initBits_4 ? 1'h0 : _GEN_2141; // @[LoadQueue.scala 308:34:@44191.4]
  assign _GEN_2143 = initBits_4 ? addrQ_4 : _GEN_2140; // @[LoadQueue.scala 308:34:@44191.4]
  assign _T_101297 = inputPriorityPorts_0_5 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44213.6]
  assign _T_101298 = inputPriorityPorts_1_5 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@44214.6]
  assign _T_101309 = _T_101297 | _T_101298; // @[LoadQueue.scala 314:26:@44219.6]
  assign _T_101310 = {_T_101298,_T_101297}; // @[OneHot.scala 18:45:@44221.8]
  assign _T_101311 = _T_101310[1]; // @[CircuitMath.scala 30:8:@44222.8]
  assign _GEN_2145 = _T_101311 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@44223.8]
  assign _GEN_2146 = _T_101309 ? _GEN_2145 : addrQ_5; // @[LoadQueue.scala 314:36:@44220.6]
  assign _GEN_2147 = _T_101309 ? 1'h1 : addrKnown_5; // @[LoadQueue.scala 314:36:@44220.6]
  assign _GEN_2148 = initBits_5 ? 1'h0 : _GEN_2147; // @[LoadQueue.scala 308:34:@44209.4]
  assign _GEN_2149 = initBits_5 ? addrQ_5 : _GEN_2146; // @[LoadQueue.scala 308:34:@44209.4]
  assign _T_101315 = inputPriorityPorts_0_6 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44231.6]
  assign _T_101316 = inputPriorityPorts_1_6 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@44232.6]
  assign _T_101327 = _T_101315 | _T_101316; // @[LoadQueue.scala 314:26:@44237.6]
  assign _T_101328 = {_T_101316,_T_101315}; // @[OneHot.scala 18:45:@44239.8]
  assign _T_101329 = _T_101328[1]; // @[CircuitMath.scala 30:8:@44240.8]
  assign _GEN_2151 = _T_101329 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@44241.8]
  assign _GEN_2152 = _T_101327 ? _GEN_2151 : addrQ_6; // @[LoadQueue.scala 314:36:@44238.6]
  assign _GEN_2153 = _T_101327 ? 1'h1 : addrKnown_6; // @[LoadQueue.scala 314:36:@44238.6]
  assign _GEN_2154 = initBits_6 ? 1'h0 : _GEN_2153; // @[LoadQueue.scala 308:34:@44227.4]
  assign _GEN_2155 = initBits_6 ? addrQ_6 : _GEN_2152; // @[LoadQueue.scala 308:34:@44227.4]
  assign _T_101333 = inputPriorityPorts_0_7 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44249.6]
  assign _T_101334 = inputPriorityPorts_1_7 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@44250.6]
  assign _T_101345 = _T_101333 | _T_101334; // @[LoadQueue.scala 314:26:@44255.6]
  assign _T_101346 = {_T_101334,_T_101333}; // @[OneHot.scala 18:45:@44257.8]
  assign _T_101347 = _T_101346[1]; // @[CircuitMath.scala 30:8:@44258.8]
  assign _GEN_2157 = _T_101347 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@44259.8]
  assign _GEN_2158 = _T_101345 ? _GEN_2157 : addrQ_7; // @[LoadQueue.scala 314:36:@44256.6]
  assign _GEN_2159 = _T_101345 ? 1'h1 : addrKnown_7; // @[LoadQueue.scala 314:36:@44256.6]
  assign _GEN_2160 = initBits_7 ? 1'h0 : _GEN_2159; // @[LoadQueue.scala 308:34:@44245.4]
  assign _GEN_2161 = initBits_7 ? addrQ_7 : _GEN_2158; // @[LoadQueue.scala 308:34:@44245.4]
  assign _T_101351 = inputPriorityPorts_0_8 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44267.6]
  assign _T_101352 = inputPriorityPorts_1_8 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@44268.6]
  assign _T_101363 = _T_101351 | _T_101352; // @[LoadQueue.scala 314:26:@44273.6]
  assign _T_101364 = {_T_101352,_T_101351}; // @[OneHot.scala 18:45:@44275.8]
  assign _T_101365 = _T_101364[1]; // @[CircuitMath.scala 30:8:@44276.8]
  assign _GEN_2163 = _T_101365 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@44277.8]
  assign _GEN_2164 = _T_101363 ? _GEN_2163 : addrQ_8; // @[LoadQueue.scala 314:36:@44274.6]
  assign _GEN_2165 = _T_101363 ? 1'h1 : addrKnown_8; // @[LoadQueue.scala 314:36:@44274.6]
  assign _GEN_2166 = initBits_8 ? 1'h0 : _GEN_2165; // @[LoadQueue.scala 308:34:@44263.4]
  assign _GEN_2167 = initBits_8 ? addrQ_8 : _GEN_2164; // @[LoadQueue.scala 308:34:@44263.4]
  assign _T_101369 = inputPriorityPorts_0_9 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44285.6]
  assign _T_101370 = inputPriorityPorts_1_9 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@44286.6]
  assign _T_101381 = _T_101369 | _T_101370; // @[LoadQueue.scala 314:26:@44291.6]
  assign _T_101382 = {_T_101370,_T_101369}; // @[OneHot.scala 18:45:@44293.8]
  assign _T_101383 = _T_101382[1]; // @[CircuitMath.scala 30:8:@44294.8]
  assign _GEN_2169 = _T_101383 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@44295.8]
  assign _GEN_2170 = _T_101381 ? _GEN_2169 : addrQ_9; // @[LoadQueue.scala 314:36:@44292.6]
  assign _GEN_2171 = _T_101381 ? 1'h1 : addrKnown_9; // @[LoadQueue.scala 314:36:@44292.6]
  assign _GEN_2172 = initBits_9 ? 1'h0 : _GEN_2171; // @[LoadQueue.scala 308:34:@44281.4]
  assign _GEN_2173 = initBits_9 ? addrQ_9 : _GEN_2170; // @[LoadQueue.scala 308:34:@44281.4]
  assign _T_101387 = inputPriorityPorts_0_10 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44303.6]
  assign _T_101388 = inputPriorityPorts_1_10 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@44304.6]
  assign _T_101399 = _T_101387 | _T_101388; // @[LoadQueue.scala 314:26:@44309.6]
  assign _T_101400 = {_T_101388,_T_101387}; // @[OneHot.scala 18:45:@44311.8]
  assign _T_101401 = _T_101400[1]; // @[CircuitMath.scala 30:8:@44312.8]
  assign _GEN_2175 = _T_101401 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@44313.8]
  assign _GEN_2176 = _T_101399 ? _GEN_2175 : addrQ_10; // @[LoadQueue.scala 314:36:@44310.6]
  assign _GEN_2177 = _T_101399 ? 1'h1 : addrKnown_10; // @[LoadQueue.scala 314:36:@44310.6]
  assign _GEN_2178 = initBits_10 ? 1'h0 : _GEN_2177; // @[LoadQueue.scala 308:34:@44299.4]
  assign _GEN_2179 = initBits_10 ? addrQ_10 : _GEN_2176; // @[LoadQueue.scala 308:34:@44299.4]
  assign _T_101405 = inputPriorityPorts_0_11 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44321.6]
  assign _T_101406 = inputPriorityPorts_1_11 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@44322.6]
  assign _T_101417 = _T_101405 | _T_101406; // @[LoadQueue.scala 314:26:@44327.6]
  assign _T_101418 = {_T_101406,_T_101405}; // @[OneHot.scala 18:45:@44329.8]
  assign _T_101419 = _T_101418[1]; // @[CircuitMath.scala 30:8:@44330.8]
  assign _GEN_2181 = _T_101419 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@44331.8]
  assign _GEN_2182 = _T_101417 ? _GEN_2181 : addrQ_11; // @[LoadQueue.scala 314:36:@44328.6]
  assign _GEN_2183 = _T_101417 ? 1'h1 : addrKnown_11; // @[LoadQueue.scala 314:36:@44328.6]
  assign _GEN_2184 = initBits_11 ? 1'h0 : _GEN_2183; // @[LoadQueue.scala 308:34:@44317.4]
  assign _GEN_2185 = initBits_11 ? addrQ_11 : _GEN_2182; // @[LoadQueue.scala 308:34:@44317.4]
  assign _T_101423 = inputPriorityPorts_0_12 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44339.6]
  assign _T_101424 = inputPriorityPorts_1_12 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@44340.6]
  assign _T_101435 = _T_101423 | _T_101424; // @[LoadQueue.scala 314:26:@44345.6]
  assign _T_101436 = {_T_101424,_T_101423}; // @[OneHot.scala 18:45:@44347.8]
  assign _T_101437 = _T_101436[1]; // @[CircuitMath.scala 30:8:@44348.8]
  assign _GEN_2187 = _T_101437 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@44349.8]
  assign _GEN_2188 = _T_101435 ? _GEN_2187 : addrQ_12; // @[LoadQueue.scala 314:36:@44346.6]
  assign _GEN_2189 = _T_101435 ? 1'h1 : addrKnown_12; // @[LoadQueue.scala 314:36:@44346.6]
  assign _GEN_2190 = initBits_12 ? 1'h0 : _GEN_2189; // @[LoadQueue.scala 308:34:@44335.4]
  assign _GEN_2191 = initBits_12 ? addrQ_12 : _GEN_2188; // @[LoadQueue.scala 308:34:@44335.4]
  assign _T_101441 = inputPriorityPorts_0_13 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44357.6]
  assign _T_101442 = inputPriorityPorts_1_13 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@44358.6]
  assign _T_101453 = _T_101441 | _T_101442; // @[LoadQueue.scala 314:26:@44363.6]
  assign _T_101454 = {_T_101442,_T_101441}; // @[OneHot.scala 18:45:@44365.8]
  assign _T_101455 = _T_101454[1]; // @[CircuitMath.scala 30:8:@44366.8]
  assign _GEN_2193 = _T_101455 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@44367.8]
  assign _GEN_2194 = _T_101453 ? _GEN_2193 : addrQ_13; // @[LoadQueue.scala 314:36:@44364.6]
  assign _GEN_2195 = _T_101453 ? 1'h1 : addrKnown_13; // @[LoadQueue.scala 314:36:@44364.6]
  assign _GEN_2196 = initBits_13 ? 1'h0 : _GEN_2195; // @[LoadQueue.scala 308:34:@44353.4]
  assign _GEN_2197 = initBits_13 ? addrQ_13 : _GEN_2194; // @[LoadQueue.scala 308:34:@44353.4]
  assign _T_101459 = inputPriorityPorts_0_14 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44375.6]
  assign _T_101460 = inputPriorityPorts_1_14 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@44376.6]
  assign _T_101471 = _T_101459 | _T_101460; // @[LoadQueue.scala 314:26:@44381.6]
  assign _T_101472 = {_T_101460,_T_101459}; // @[OneHot.scala 18:45:@44383.8]
  assign _T_101473 = _T_101472[1]; // @[CircuitMath.scala 30:8:@44384.8]
  assign _GEN_2199 = _T_101473 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@44385.8]
  assign _GEN_2200 = _T_101471 ? _GEN_2199 : addrQ_14; // @[LoadQueue.scala 314:36:@44382.6]
  assign _GEN_2201 = _T_101471 ? 1'h1 : addrKnown_14; // @[LoadQueue.scala 314:36:@44382.6]
  assign _GEN_2202 = initBits_14 ? 1'h0 : _GEN_2201; // @[LoadQueue.scala 308:34:@44371.4]
  assign _GEN_2203 = initBits_14 ? addrQ_14 : _GEN_2200; // @[LoadQueue.scala 308:34:@44371.4]
  assign _T_101477 = inputPriorityPorts_0_15 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44393.6]
  assign _T_101478 = inputPriorityPorts_1_15 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@44394.6]
  assign _T_101489 = _T_101477 | _T_101478; // @[LoadQueue.scala 314:26:@44399.6]
  assign _T_101490 = {_T_101478,_T_101477}; // @[OneHot.scala 18:45:@44401.8]
  assign _T_101491 = _T_101490[1]; // @[CircuitMath.scala 30:8:@44402.8]
  assign _GEN_2205 = _T_101491 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@44403.8]
  assign _GEN_2206 = _T_101489 ? _GEN_2205 : addrQ_15; // @[LoadQueue.scala 314:36:@44400.6]
  assign _GEN_2207 = _T_101489 ? 1'h1 : addrKnown_15; // @[LoadQueue.scala 314:36:@44400.6]
  assign _GEN_2208 = initBits_15 ? 1'h0 : _GEN_2207; // @[LoadQueue.scala 308:34:@44389.4]
  assign _GEN_2209 = initBits_15 ? addrQ_15 : _GEN_2206; // @[LoadQueue.scala 308:34:@44389.4]
  assign _T_101515 = outputPriorityPorts_0_0 & dataKnown_0; // @[LoadQueue.scala 326:108:@44408.4]
  assign _T_101517 = loadCompleted_0 == 1'h0; // @[LoadQueue.scala 327:34:@44409.4]
  assign _T_101518 = _T_101515 & _T_101517; // @[LoadQueue.scala 327:31:@44410.4]
  assign _T_101519 = _T_101518 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44411.4]
  assign _T_101520 = outputPriorityPorts_1_0 & dataKnown_0; // @[LoadQueue.scala 326:108:@44412.4]
  assign _T_101523 = _T_101520 & _T_101517; // @[LoadQueue.scala 327:31:@44414.4]
  assign _T_101524 = _T_101523 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@44415.4]
  assign loadCompleting_0 = _T_101519 | _T_101524; // @[LoadQueue.scala 328:51:@44420.4]
  assign _T_101536 = outputPriorityPorts_0_1 & dataKnown_1; // @[LoadQueue.scala 326:108:@44422.4]
  assign _T_101538 = loadCompleted_1 == 1'h0; // @[LoadQueue.scala 327:34:@44423.4]
  assign _T_101539 = _T_101536 & _T_101538; // @[LoadQueue.scala 327:31:@44424.4]
  assign _T_101540 = _T_101539 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44425.4]
  assign _T_101541 = outputPriorityPorts_1_1 & dataKnown_1; // @[LoadQueue.scala 326:108:@44426.4]
  assign _T_101544 = _T_101541 & _T_101538; // @[LoadQueue.scala 327:31:@44428.4]
  assign _T_101545 = _T_101544 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@44429.4]
  assign loadCompleting_1 = _T_101540 | _T_101545; // @[LoadQueue.scala 328:51:@44434.4]
  assign _T_101557 = outputPriorityPorts_0_2 & dataKnown_2; // @[LoadQueue.scala 326:108:@44436.4]
  assign _T_101559 = loadCompleted_2 == 1'h0; // @[LoadQueue.scala 327:34:@44437.4]
  assign _T_101560 = _T_101557 & _T_101559; // @[LoadQueue.scala 327:31:@44438.4]
  assign _T_101561 = _T_101560 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44439.4]
  assign _T_101562 = outputPriorityPorts_1_2 & dataKnown_2; // @[LoadQueue.scala 326:108:@44440.4]
  assign _T_101565 = _T_101562 & _T_101559; // @[LoadQueue.scala 327:31:@44442.4]
  assign _T_101566 = _T_101565 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@44443.4]
  assign loadCompleting_2 = _T_101561 | _T_101566; // @[LoadQueue.scala 328:51:@44448.4]
  assign _T_101578 = outputPriorityPorts_0_3 & dataKnown_3; // @[LoadQueue.scala 326:108:@44450.4]
  assign _T_101580 = loadCompleted_3 == 1'h0; // @[LoadQueue.scala 327:34:@44451.4]
  assign _T_101581 = _T_101578 & _T_101580; // @[LoadQueue.scala 327:31:@44452.4]
  assign _T_101582 = _T_101581 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44453.4]
  assign _T_101583 = outputPriorityPorts_1_3 & dataKnown_3; // @[LoadQueue.scala 326:108:@44454.4]
  assign _T_101586 = _T_101583 & _T_101580; // @[LoadQueue.scala 327:31:@44456.4]
  assign _T_101587 = _T_101586 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@44457.4]
  assign loadCompleting_3 = _T_101582 | _T_101587; // @[LoadQueue.scala 328:51:@44462.4]
  assign _T_101599 = outputPriorityPorts_0_4 & dataKnown_4; // @[LoadQueue.scala 326:108:@44464.4]
  assign _T_101601 = loadCompleted_4 == 1'h0; // @[LoadQueue.scala 327:34:@44465.4]
  assign _T_101602 = _T_101599 & _T_101601; // @[LoadQueue.scala 327:31:@44466.4]
  assign _T_101603 = _T_101602 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44467.4]
  assign _T_101604 = outputPriorityPorts_1_4 & dataKnown_4; // @[LoadQueue.scala 326:108:@44468.4]
  assign _T_101607 = _T_101604 & _T_101601; // @[LoadQueue.scala 327:31:@44470.4]
  assign _T_101608 = _T_101607 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@44471.4]
  assign loadCompleting_4 = _T_101603 | _T_101608; // @[LoadQueue.scala 328:51:@44476.4]
  assign _T_101620 = outputPriorityPorts_0_5 & dataKnown_5; // @[LoadQueue.scala 326:108:@44478.4]
  assign _T_101622 = loadCompleted_5 == 1'h0; // @[LoadQueue.scala 327:34:@44479.4]
  assign _T_101623 = _T_101620 & _T_101622; // @[LoadQueue.scala 327:31:@44480.4]
  assign _T_101624 = _T_101623 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44481.4]
  assign _T_101625 = outputPriorityPorts_1_5 & dataKnown_5; // @[LoadQueue.scala 326:108:@44482.4]
  assign _T_101628 = _T_101625 & _T_101622; // @[LoadQueue.scala 327:31:@44484.4]
  assign _T_101629 = _T_101628 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@44485.4]
  assign loadCompleting_5 = _T_101624 | _T_101629; // @[LoadQueue.scala 328:51:@44490.4]
  assign _T_101641 = outputPriorityPorts_0_6 & dataKnown_6; // @[LoadQueue.scala 326:108:@44492.4]
  assign _T_101643 = loadCompleted_6 == 1'h0; // @[LoadQueue.scala 327:34:@44493.4]
  assign _T_101644 = _T_101641 & _T_101643; // @[LoadQueue.scala 327:31:@44494.4]
  assign _T_101645 = _T_101644 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44495.4]
  assign _T_101646 = outputPriorityPorts_1_6 & dataKnown_6; // @[LoadQueue.scala 326:108:@44496.4]
  assign _T_101649 = _T_101646 & _T_101643; // @[LoadQueue.scala 327:31:@44498.4]
  assign _T_101650 = _T_101649 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@44499.4]
  assign loadCompleting_6 = _T_101645 | _T_101650; // @[LoadQueue.scala 328:51:@44504.4]
  assign _T_101662 = outputPriorityPorts_0_7 & dataKnown_7; // @[LoadQueue.scala 326:108:@44506.4]
  assign _T_101664 = loadCompleted_7 == 1'h0; // @[LoadQueue.scala 327:34:@44507.4]
  assign _T_101665 = _T_101662 & _T_101664; // @[LoadQueue.scala 327:31:@44508.4]
  assign _T_101666 = _T_101665 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44509.4]
  assign _T_101667 = outputPriorityPorts_1_7 & dataKnown_7; // @[LoadQueue.scala 326:108:@44510.4]
  assign _T_101670 = _T_101667 & _T_101664; // @[LoadQueue.scala 327:31:@44512.4]
  assign _T_101671 = _T_101670 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@44513.4]
  assign loadCompleting_7 = _T_101666 | _T_101671; // @[LoadQueue.scala 328:51:@44518.4]
  assign _T_101683 = outputPriorityPorts_0_8 & dataKnown_8; // @[LoadQueue.scala 326:108:@44520.4]
  assign _T_101685 = loadCompleted_8 == 1'h0; // @[LoadQueue.scala 327:34:@44521.4]
  assign _T_101686 = _T_101683 & _T_101685; // @[LoadQueue.scala 327:31:@44522.4]
  assign _T_101687 = _T_101686 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44523.4]
  assign _T_101688 = outputPriorityPorts_1_8 & dataKnown_8; // @[LoadQueue.scala 326:108:@44524.4]
  assign _T_101691 = _T_101688 & _T_101685; // @[LoadQueue.scala 327:31:@44526.4]
  assign _T_101692 = _T_101691 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@44527.4]
  assign loadCompleting_8 = _T_101687 | _T_101692; // @[LoadQueue.scala 328:51:@44532.4]
  assign _T_101704 = outputPriorityPorts_0_9 & dataKnown_9; // @[LoadQueue.scala 326:108:@44534.4]
  assign _T_101706 = loadCompleted_9 == 1'h0; // @[LoadQueue.scala 327:34:@44535.4]
  assign _T_101707 = _T_101704 & _T_101706; // @[LoadQueue.scala 327:31:@44536.4]
  assign _T_101708 = _T_101707 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44537.4]
  assign _T_101709 = outputPriorityPorts_1_9 & dataKnown_9; // @[LoadQueue.scala 326:108:@44538.4]
  assign _T_101712 = _T_101709 & _T_101706; // @[LoadQueue.scala 327:31:@44540.4]
  assign _T_101713 = _T_101712 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@44541.4]
  assign loadCompleting_9 = _T_101708 | _T_101713; // @[LoadQueue.scala 328:51:@44546.4]
  assign _T_101725 = outputPriorityPorts_0_10 & dataKnown_10; // @[LoadQueue.scala 326:108:@44548.4]
  assign _T_101727 = loadCompleted_10 == 1'h0; // @[LoadQueue.scala 327:34:@44549.4]
  assign _T_101728 = _T_101725 & _T_101727; // @[LoadQueue.scala 327:31:@44550.4]
  assign _T_101729 = _T_101728 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44551.4]
  assign _T_101730 = outputPriorityPorts_1_10 & dataKnown_10; // @[LoadQueue.scala 326:108:@44552.4]
  assign _T_101733 = _T_101730 & _T_101727; // @[LoadQueue.scala 327:31:@44554.4]
  assign _T_101734 = _T_101733 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@44555.4]
  assign loadCompleting_10 = _T_101729 | _T_101734; // @[LoadQueue.scala 328:51:@44560.4]
  assign _T_101746 = outputPriorityPorts_0_11 & dataKnown_11; // @[LoadQueue.scala 326:108:@44562.4]
  assign _T_101748 = loadCompleted_11 == 1'h0; // @[LoadQueue.scala 327:34:@44563.4]
  assign _T_101749 = _T_101746 & _T_101748; // @[LoadQueue.scala 327:31:@44564.4]
  assign _T_101750 = _T_101749 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44565.4]
  assign _T_101751 = outputPriorityPorts_1_11 & dataKnown_11; // @[LoadQueue.scala 326:108:@44566.4]
  assign _T_101754 = _T_101751 & _T_101748; // @[LoadQueue.scala 327:31:@44568.4]
  assign _T_101755 = _T_101754 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@44569.4]
  assign loadCompleting_11 = _T_101750 | _T_101755; // @[LoadQueue.scala 328:51:@44574.4]
  assign _T_101767 = outputPriorityPorts_0_12 & dataKnown_12; // @[LoadQueue.scala 326:108:@44576.4]
  assign _T_101769 = loadCompleted_12 == 1'h0; // @[LoadQueue.scala 327:34:@44577.4]
  assign _T_101770 = _T_101767 & _T_101769; // @[LoadQueue.scala 327:31:@44578.4]
  assign _T_101771 = _T_101770 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44579.4]
  assign _T_101772 = outputPriorityPorts_1_12 & dataKnown_12; // @[LoadQueue.scala 326:108:@44580.4]
  assign _T_101775 = _T_101772 & _T_101769; // @[LoadQueue.scala 327:31:@44582.4]
  assign _T_101776 = _T_101775 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@44583.4]
  assign loadCompleting_12 = _T_101771 | _T_101776; // @[LoadQueue.scala 328:51:@44588.4]
  assign _T_101788 = outputPriorityPorts_0_13 & dataKnown_13; // @[LoadQueue.scala 326:108:@44590.4]
  assign _T_101790 = loadCompleted_13 == 1'h0; // @[LoadQueue.scala 327:34:@44591.4]
  assign _T_101791 = _T_101788 & _T_101790; // @[LoadQueue.scala 327:31:@44592.4]
  assign _T_101792 = _T_101791 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44593.4]
  assign _T_101793 = outputPriorityPorts_1_13 & dataKnown_13; // @[LoadQueue.scala 326:108:@44594.4]
  assign _T_101796 = _T_101793 & _T_101790; // @[LoadQueue.scala 327:31:@44596.4]
  assign _T_101797 = _T_101796 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@44597.4]
  assign loadCompleting_13 = _T_101792 | _T_101797; // @[LoadQueue.scala 328:51:@44602.4]
  assign _T_101809 = outputPriorityPorts_0_14 & dataKnown_14; // @[LoadQueue.scala 326:108:@44604.4]
  assign _T_101811 = loadCompleted_14 == 1'h0; // @[LoadQueue.scala 327:34:@44605.4]
  assign _T_101812 = _T_101809 & _T_101811; // @[LoadQueue.scala 327:31:@44606.4]
  assign _T_101813 = _T_101812 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44607.4]
  assign _T_101814 = outputPriorityPorts_1_14 & dataKnown_14; // @[LoadQueue.scala 326:108:@44608.4]
  assign _T_101817 = _T_101814 & _T_101811; // @[LoadQueue.scala 327:31:@44610.4]
  assign _T_101818 = _T_101817 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@44611.4]
  assign loadCompleting_14 = _T_101813 | _T_101818; // @[LoadQueue.scala 328:51:@44616.4]
  assign _T_101830 = outputPriorityPorts_0_15 & dataKnown_15; // @[LoadQueue.scala 326:108:@44618.4]
  assign _T_101832 = loadCompleted_15 == 1'h0; // @[LoadQueue.scala 327:34:@44619.4]
  assign _T_101833 = _T_101830 & _T_101832; // @[LoadQueue.scala 327:31:@44620.4]
  assign _T_101834 = _T_101833 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44621.4]
  assign _T_101835 = outputPriorityPorts_1_15 & dataKnown_15; // @[LoadQueue.scala 326:108:@44622.4]
  assign _T_101838 = _T_101835 & _T_101832; // @[LoadQueue.scala 327:31:@44624.4]
  assign _T_101839 = _T_101838 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@44625.4]
  assign loadCompleting_15 = _T_101834 | _T_101839; // @[LoadQueue.scala 328:51:@44630.4]
  assign _GEN_2210 = loadCompleting_0 ? 1'h1 : loadCompleted_0; // @[LoadQueue.scala 337:46:@44636.6]
  assign _GEN_2211 = initBits_0 ? 1'h0 : _GEN_2210; // @[LoadQueue.scala 335:34:@44632.4]
  assign _GEN_2212 = loadCompleting_1 ? 1'h1 : loadCompleted_1; // @[LoadQueue.scala 337:46:@44643.6]
  assign _GEN_2213 = initBits_1 ? 1'h0 : _GEN_2212; // @[LoadQueue.scala 335:34:@44639.4]
  assign _GEN_2214 = loadCompleting_2 ? 1'h1 : loadCompleted_2; // @[LoadQueue.scala 337:46:@44650.6]
  assign _GEN_2215 = initBits_2 ? 1'h0 : _GEN_2214; // @[LoadQueue.scala 335:34:@44646.4]
  assign _GEN_2216 = loadCompleting_3 ? 1'h1 : loadCompleted_3; // @[LoadQueue.scala 337:46:@44657.6]
  assign _GEN_2217 = initBits_3 ? 1'h0 : _GEN_2216; // @[LoadQueue.scala 335:34:@44653.4]
  assign _GEN_2218 = loadCompleting_4 ? 1'h1 : loadCompleted_4; // @[LoadQueue.scala 337:46:@44664.6]
  assign _GEN_2219 = initBits_4 ? 1'h0 : _GEN_2218; // @[LoadQueue.scala 335:34:@44660.4]
  assign _GEN_2220 = loadCompleting_5 ? 1'h1 : loadCompleted_5; // @[LoadQueue.scala 337:46:@44671.6]
  assign _GEN_2221 = initBits_5 ? 1'h0 : _GEN_2220; // @[LoadQueue.scala 335:34:@44667.4]
  assign _GEN_2222 = loadCompleting_6 ? 1'h1 : loadCompleted_6; // @[LoadQueue.scala 337:46:@44678.6]
  assign _GEN_2223 = initBits_6 ? 1'h0 : _GEN_2222; // @[LoadQueue.scala 335:34:@44674.4]
  assign _GEN_2224 = loadCompleting_7 ? 1'h1 : loadCompleted_7; // @[LoadQueue.scala 337:46:@44685.6]
  assign _GEN_2225 = initBits_7 ? 1'h0 : _GEN_2224; // @[LoadQueue.scala 335:34:@44681.4]
  assign _GEN_2226 = loadCompleting_8 ? 1'h1 : loadCompleted_8; // @[LoadQueue.scala 337:46:@44692.6]
  assign _GEN_2227 = initBits_8 ? 1'h0 : _GEN_2226; // @[LoadQueue.scala 335:34:@44688.4]
  assign _GEN_2228 = loadCompleting_9 ? 1'h1 : loadCompleted_9; // @[LoadQueue.scala 337:46:@44699.6]
  assign _GEN_2229 = initBits_9 ? 1'h0 : _GEN_2228; // @[LoadQueue.scala 335:34:@44695.4]
  assign _GEN_2230 = loadCompleting_10 ? 1'h1 : loadCompleted_10; // @[LoadQueue.scala 337:46:@44706.6]
  assign _GEN_2231 = initBits_10 ? 1'h0 : _GEN_2230; // @[LoadQueue.scala 335:34:@44702.4]
  assign _GEN_2232 = loadCompleting_11 ? 1'h1 : loadCompleted_11; // @[LoadQueue.scala 337:46:@44713.6]
  assign _GEN_2233 = initBits_11 ? 1'h0 : _GEN_2232; // @[LoadQueue.scala 335:34:@44709.4]
  assign _GEN_2234 = loadCompleting_12 ? 1'h1 : loadCompleted_12; // @[LoadQueue.scala 337:46:@44720.6]
  assign _GEN_2235 = initBits_12 ? 1'h0 : _GEN_2234; // @[LoadQueue.scala 335:34:@44716.4]
  assign _GEN_2236 = loadCompleting_13 ? 1'h1 : loadCompleted_13; // @[LoadQueue.scala 337:46:@44727.6]
  assign _GEN_2237 = initBits_13 ? 1'h0 : _GEN_2236; // @[LoadQueue.scala 335:34:@44723.4]
  assign _GEN_2238 = loadCompleting_14 ? 1'h1 : loadCompleted_14; // @[LoadQueue.scala 337:46:@44734.6]
  assign _GEN_2239 = initBits_14 ? 1'h0 : _GEN_2238; // @[LoadQueue.scala 335:34:@44730.4]
  assign _GEN_2240 = loadCompleting_15 ? 1'h1 : loadCompleted_15; // @[LoadQueue.scala 337:46:@44741.6]
  assign _GEN_2241 = initBits_15 ? 1'h0 : _GEN_2240; // @[LoadQueue.scala 335:34:@44737.4]
  assign _T_101971 = _T_101518 | _T_101539; // @[LoadQueue.scala 348:24:@44810.4]
  assign _T_101972 = _T_101971 | _T_101560; // @[LoadQueue.scala 348:24:@44811.4]
  assign _T_101973 = _T_101972 | _T_101581; // @[LoadQueue.scala 348:24:@44812.4]
  assign _T_101974 = _T_101973 | _T_101602; // @[LoadQueue.scala 348:24:@44813.4]
  assign _T_101975 = _T_101974 | _T_101623; // @[LoadQueue.scala 348:24:@44814.4]
  assign _T_101976 = _T_101975 | _T_101644; // @[LoadQueue.scala 348:24:@44815.4]
  assign _T_101977 = _T_101976 | _T_101665; // @[LoadQueue.scala 348:24:@44816.4]
  assign _T_101978 = _T_101977 | _T_101686; // @[LoadQueue.scala 348:24:@44817.4]
  assign _T_101979 = _T_101978 | _T_101707; // @[LoadQueue.scala 348:24:@44818.4]
  assign _T_101980 = _T_101979 | _T_101728; // @[LoadQueue.scala 348:24:@44819.4]
  assign _T_101981 = _T_101980 | _T_101749; // @[LoadQueue.scala 348:24:@44820.4]
  assign _T_101982 = _T_101981 | _T_101770; // @[LoadQueue.scala 348:24:@44821.4]
  assign _T_101983 = _T_101982 | _T_101791; // @[LoadQueue.scala 348:24:@44822.4]
  assign _T_101984 = _T_101983 | _T_101812; // @[LoadQueue.scala 348:24:@44823.4]
  assign _T_101985 = _T_101984 | _T_101833; // @[LoadQueue.scala 348:24:@44824.4]
  assign _T_102002 = _T_101812 ? 4'he : 4'hf; // @[Mux.scala 31:69:@44826.6]
  assign _T_102003 = _T_101791 ? 4'hd : _T_102002; // @[Mux.scala 31:69:@44827.6]
  assign _T_102004 = _T_101770 ? 4'hc : _T_102003; // @[Mux.scala 31:69:@44828.6]
  assign _T_102005 = _T_101749 ? 4'hb : _T_102004; // @[Mux.scala 31:69:@44829.6]
  assign _T_102006 = _T_101728 ? 4'ha : _T_102005; // @[Mux.scala 31:69:@44830.6]
  assign _T_102007 = _T_101707 ? 4'h9 : _T_102006; // @[Mux.scala 31:69:@44831.6]
  assign _T_102008 = _T_101686 ? 4'h8 : _T_102007; // @[Mux.scala 31:69:@44832.6]
  assign _T_102009 = _T_101665 ? 4'h7 : _T_102008; // @[Mux.scala 31:69:@44833.6]
  assign _T_102010 = _T_101644 ? 4'h6 : _T_102009; // @[Mux.scala 31:69:@44834.6]
  assign _T_102011 = _T_101623 ? 4'h5 : _T_102010; // @[Mux.scala 31:69:@44835.6]
  assign _T_102012 = _T_101602 ? 4'h4 : _T_102011; // @[Mux.scala 31:69:@44836.6]
  assign _T_102013 = _T_101581 ? 4'h3 : _T_102012; // @[Mux.scala 31:69:@44837.6]
  assign _T_102014 = _T_101560 ? 4'h2 : _T_102013; // @[Mux.scala 31:69:@44838.6]
  assign _T_102015 = _T_101539 ? 4'h1 : _T_102014; // @[Mux.scala 31:69:@44839.6]
  assign _T_102016 = _T_101518 ? 4'h0 : _T_102015; // @[Mux.scala 31:69:@44840.6]
  assign _GEN_2243 = 4'h1 == _T_102016 ? dataQ_1 : dataQ_0; // @[LoadQueue.scala 349:37:@44841.6]
  assign _GEN_2244 = 4'h2 == _T_102016 ? dataQ_2 : _GEN_2243; // @[LoadQueue.scala 349:37:@44841.6]
  assign _GEN_2245 = 4'h3 == _T_102016 ? dataQ_3 : _GEN_2244; // @[LoadQueue.scala 349:37:@44841.6]
  assign _GEN_2246 = 4'h4 == _T_102016 ? dataQ_4 : _GEN_2245; // @[LoadQueue.scala 349:37:@44841.6]
  assign _GEN_2247 = 4'h5 == _T_102016 ? dataQ_5 : _GEN_2246; // @[LoadQueue.scala 349:37:@44841.6]
  assign _GEN_2248 = 4'h6 == _T_102016 ? dataQ_6 : _GEN_2247; // @[LoadQueue.scala 349:37:@44841.6]
  assign _GEN_2249 = 4'h7 == _T_102016 ? dataQ_7 : _GEN_2248; // @[LoadQueue.scala 349:37:@44841.6]
  assign _GEN_2250 = 4'h8 == _T_102016 ? dataQ_8 : _GEN_2249; // @[LoadQueue.scala 349:37:@44841.6]
  assign _GEN_2251 = 4'h9 == _T_102016 ? dataQ_9 : _GEN_2250; // @[LoadQueue.scala 349:37:@44841.6]
  assign _GEN_2252 = 4'ha == _T_102016 ? dataQ_10 : _GEN_2251; // @[LoadQueue.scala 349:37:@44841.6]
  assign _GEN_2253 = 4'hb == _T_102016 ? dataQ_11 : _GEN_2252; // @[LoadQueue.scala 349:37:@44841.6]
  assign _GEN_2254 = 4'hc == _T_102016 ? dataQ_12 : _GEN_2253; // @[LoadQueue.scala 349:37:@44841.6]
  assign _GEN_2255 = 4'hd == _T_102016 ? dataQ_13 : _GEN_2254; // @[LoadQueue.scala 349:37:@44841.6]
  assign _GEN_2256 = 4'he == _T_102016 ? dataQ_14 : _GEN_2255; // @[LoadQueue.scala 349:37:@44841.6]
  assign _GEN_2257 = 4'hf == _T_102016 ? dataQ_15 : _GEN_2256; // @[LoadQueue.scala 349:37:@44841.6]
  assign _T_102111 = _T_101523 | _T_101544; // @[LoadQueue.scala 348:24:@44914.4]
  assign _T_102112 = _T_102111 | _T_101565; // @[LoadQueue.scala 348:24:@44915.4]
  assign _T_102113 = _T_102112 | _T_101586; // @[LoadQueue.scala 348:24:@44916.4]
  assign _T_102114 = _T_102113 | _T_101607; // @[LoadQueue.scala 348:24:@44917.4]
  assign _T_102115 = _T_102114 | _T_101628; // @[LoadQueue.scala 348:24:@44918.4]
  assign _T_102116 = _T_102115 | _T_101649; // @[LoadQueue.scala 348:24:@44919.4]
  assign _T_102117 = _T_102116 | _T_101670; // @[LoadQueue.scala 348:24:@44920.4]
  assign _T_102118 = _T_102117 | _T_101691; // @[LoadQueue.scala 348:24:@44921.4]
  assign _T_102119 = _T_102118 | _T_101712; // @[LoadQueue.scala 348:24:@44922.4]
  assign _T_102120 = _T_102119 | _T_101733; // @[LoadQueue.scala 348:24:@44923.4]
  assign _T_102121 = _T_102120 | _T_101754; // @[LoadQueue.scala 348:24:@44924.4]
  assign _T_102122 = _T_102121 | _T_101775; // @[LoadQueue.scala 348:24:@44925.4]
  assign _T_102123 = _T_102122 | _T_101796; // @[LoadQueue.scala 348:24:@44926.4]
  assign _T_102124 = _T_102123 | _T_101817; // @[LoadQueue.scala 348:24:@44927.4]
  assign _T_102125 = _T_102124 | _T_101838; // @[LoadQueue.scala 348:24:@44928.4]
  assign _T_102142 = _T_101817 ? 4'he : 4'hf; // @[Mux.scala 31:69:@44930.6]
  assign _T_102143 = _T_101796 ? 4'hd : _T_102142; // @[Mux.scala 31:69:@44931.6]
  assign _T_102144 = _T_101775 ? 4'hc : _T_102143; // @[Mux.scala 31:69:@44932.6]
  assign _T_102145 = _T_101754 ? 4'hb : _T_102144; // @[Mux.scala 31:69:@44933.6]
  assign _T_102146 = _T_101733 ? 4'ha : _T_102145; // @[Mux.scala 31:69:@44934.6]
  assign _T_102147 = _T_101712 ? 4'h9 : _T_102146; // @[Mux.scala 31:69:@44935.6]
  assign _T_102148 = _T_101691 ? 4'h8 : _T_102147; // @[Mux.scala 31:69:@44936.6]
  assign _T_102149 = _T_101670 ? 4'h7 : _T_102148; // @[Mux.scala 31:69:@44937.6]
  assign _T_102150 = _T_101649 ? 4'h6 : _T_102149; // @[Mux.scala 31:69:@44938.6]
  assign _T_102151 = _T_101628 ? 4'h5 : _T_102150; // @[Mux.scala 31:69:@44939.6]
  assign _T_102152 = _T_101607 ? 4'h4 : _T_102151; // @[Mux.scala 31:69:@44940.6]
  assign _T_102153 = _T_101586 ? 4'h3 : _T_102152; // @[Mux.scala 31:69:@44941.6]
  assign _T_102154 = _T_101565 ? 4'h2 : _T_102153; // @[Mux.scala 31:69:@44942.6]
  assign _T_102155 = _T_101544 ? 4'h1 : _T_102154; // @[Mux.scala 31:69:@44943.6]
  assign _T_102156 = _T_101523 ? 4'h0 : _T_102155; // @[Mux.scala 31:69:@44944.6]
  assign _GEN_2261 = 4'h1 == _T_102156 ? dataQ_1 : dataQ_0; // @[LoadQueue.scala 349:37:@44945.6]
  assign _GEN_2262 = 4'h2 == _T_102156 ? dataQ_2 : _GEN_2261; // @[LoadQueue.scala 349:37:@44945.6]
  assign _GEN_2263 = 4'h3 == _T_102156 ? dataQ_3 : _GEN_2262; // @[LoadQueue.scala 349:37:@44945.6]
  assign _GEN_2264 = 4'h4 == _T_102156 ? dataQ_4 : _GEN_2263; // @[LoadQueue.scala 349:37:@44945.6]
  assign _GEN_2265 = 4'h5 == _T_102156 ? dataQ_5 : _GEN_2264; // @[LoadQueue.scala 349:37:@44945.6]
  assign _GEN_2266 = 4'h6 == _T_102156 ? dataQ_6 : _GEN_2265; // @[LoadQueue.scala 349:37:@44945.6]
  assign _GEN_2267 = 4'h7 == _T_102156 ? dataQ_7 : _GEN_2266; // @[LoadQueue.scala 349:37:@44945.6]
  assign _GEN_2268 = 4'h8 == _T_102156 ? dataQ_8 : _GEN_2267; // @[LoadQueue.scala 349:37:@44945.6]
  assign _GEN_2269 = 4'h9 == _T_102156 ? dataQ_9 : _GEN_2268; // @[LoadQueue.scala 349:37:@44945.6]
  assign _GEN_2270 = 4'ha == _T_102156 ? dataQ_10 : _GEN_2269; // @[LoadQueue.scala 349:37:@44945.6]
  assign _GEN_2271 = 4'hb == _T_102156 ? dataQ_11 : _GEN_2270; // @[LoadQueue.scala 349:37:@44945.6]
  assign _GEN_2272 = 4'hc == _T_102156 ? dataQ_12 : _GEN_2271; // @[LoadQueue.scala 349:37:@44945.6]
  assign _GEN_2273 = 4'hd == _T_102156 ? dataQ_13 : _GEN_2272; // @[LoadQueue.scala 349:37:@44945.6]
  assign _GEN_2274 = 4'he == _T_102156 ? dataQ_14 : _GEN_2273; // @[LoadQueue.scala 349:37:@44945.6]
  assign _GEN_2275 = 4'hf == _T_102156 ? dataQ_15 : _GEN_2274; // @[LoadQueue.scala 349:37:@44945.6]
  assign _GEN_2279 = 4'h1 == head ? loadCompleted_1 : loadCompleted_0; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2280 = 4'h2 == head ? loadCompleted_2 : _GEN_2279; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2281 = 4'h3 == head ? loadCompleted_3 : _GEN_2280; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2282 = 4'h4 == head ? loadCompleted_4 : _GEN_2281; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2283 = 4'h5 == head ? loadCompleted_5 : _GEN_2282; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2284 = 4'h6 == head ? loadCompleted_6 : _GEN_2283; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2285 = 4'h7 == head ? loadCompleted_7 : _GEN_2284; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2286 = 4'h8 == head ? loadCompleted_8 : _GEN_2285; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2287 = 4'h9 == head ? loadCompleted_9 : _GEN_2286; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2288 = 4'ha == head ? loadCompleted_10 : _GEN_2287; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2289 = 4'hb == head ? loadCompleted_11 : _GEN_2288; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2290 = 4'hc == head ? loadCompleted_12 : _GEN_2289; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2291 = 4'hd == head ? loadCompleted_13 : _GEN_2290; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2292 = 4'he == head ? loadCompleted_14 : _GEN_2291; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2293 = 4'hf == head ? loadCompleted_15 : _GEN_2292; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2295 = 4'h1 == head ? loadCompleting_1 : loadCompleting_0; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2296 = 4'h2 == head ? loadCompleting_2 : _GEN_2295; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2297 = 4'h3 == head ? loadCompleting_3 : _GEN_2296; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2298 = 4'h4 == head ? loadCompleting_4 : _GEN_2297; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2299 = 4'h5 == head ? loadCompleting_5 : _GEN_2298; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2300 = 4'h6 == head ? loadCompleting_6 : _GEN_2299; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2301 = 4'h7 == head ? loadCompleting_7 : _GEN_2300; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2302 = 4'h8 == head ? loadCompleting_8 : _GEN_2301; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2303 = 4'h9 == head ? loadCompleting_9 : _GEN_2302; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2304 = 4'ha == head ? loadCompleting_10 : _GEN_2303; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2305 = 4'hb == head ? loadCompleting_11 : _GEN_2304; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2306 = 4'hc == head ? loadCompleting_12 : _GEN_2305; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2307 = 4'hd == head ? loadCompleting_13 : _GEN_2306; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2308 = 4'he == head ? loadCompleting_14 : _GEN_2307; // @[LoadQueue.scala 363:29:@44952.4]
  assign _GEN_2309 = 4'hf == head ? loadCompleting_15 : _GEN_2308; // @[LoadQueue.scala 363:29:@44952.4]
  assign _T_102167 = _GEN_2293 | _GEN_2309; // @[LoadQueue.scala 363:29:@44952.4]
  assign _T_102168 = head != tail; // @[LoadQueue.scala 363:63:@44953.4]
  assign _T_102170 = io_loadEmpty == 1'h0; // @[LoadQueue.scala 363:75:@44954.4]
  assign _T_102171 = _T_102168 | _T_102170; // @[LoadQueue.scala 363:72:@44955.4]
  assign _T_102172 = _T_102167 & _T_102171; // @[LoadQueue.scala 363:54:@44956.4]
  assign _T_102175 = head + 4'h1; // @[util.scala 10:8:@44958.6]
  assign _GEN_544 = _T_102175 % 5'h10; // @[util.scala 10:14:@44959.6]
  assign _T_102176 = _GEN_544[4:0]; // @[util.scala 10:14:@44959.6]
  assign _GEN_2310 = _T_102172 ? _T_102176 : {{1'd0}, head}; // @[LoadQueue.scala 363:91:@44957.4]
  assign _GEN_2408 = {{2'd0}, io_bbNumLoads}; // @[util.scala 10:8:@44963.6]
  assign _T_102178 = tail + _GEN_2408; // @[util.scala 10:8:@44963.6]
  assign _GEN_545 = _T_102178 % 5'h10; // @[util.scala 10:14:@44964.6]
  assign _T_102179 = _GEN_545[4:0]; // @[util.scala 10:14:@44964.6]
  assign _GEN_2311 = io_bbStart ? _T_102179 : {{1'd0}, tail}; // @[LoadQueue.scala 367:20:@44962.4]
  assign _T_102181 = allocatedEntries_0 == 1'h0; // @[LoadQueue.scala 371:82:@44967.4]
  assign _T_102182 = loadCompleted_0 | _T_102181; // @[LoadQueue.scala 371:79:@44968.4]
  assign _T_102184 = allocatedEntries_1 == 1'h0; // @[LoadQueue.scala 371:82:@44969.4]
  assign _T_102185 = loadCompleted_1 | _T_102184; // @[LoadQueue.scala 371:79:@44970.4]
  assign _T_102187 = allocatedEntries_2 == 1'h0; // @[LoadQueue.scala 371:82:@44971.4]
  assign _T_102188 = loadCompleted_2 | _T_102187; // @[LoadQueue.scala 371:79:@44972.4]
  assign _T_102190 = allocatedEntries_3 == 1'h0; // @[LoadQueue.scala 371:82:@44973.4]
  assign _T_102191 = loadCompleted_3 | _T_102190; // @[LoadQueue.scala 371:79:@44974.4]
  assign _T_102193 = allocatedEntries_4 == 1'h0; // @[LoadQueue.scala 371:82:@44975.4]
  assign _T_102194 = loadCompleted_4 | _T_102193; // @[LoadQueue.scala 371:79:@44976.4]
  assign _T_102196 = allocatedEntries_5 == 1'h0; // @[LoadQueue.scala 371:82:@44977.4]
  assign _T_102197 = loadCompleted_5 | _T_102196; // @[LoadQueue.scala 371:79:@44978.4]
  assign _T_102199 = allocatedEntries_6 == 1'h0; // @[LoadQueue.scala 371:82:@44979.4]
  assign _T_102200 = loadCompleted_6 | _T_102199; // @[LoadQueue.scala 371:79:@44980.4]
  assign _T_102202 = allocatedEntries_7 == 1'h0; // @[LoadQueue.scala 371:82:@44981.4]
  assign _T_102203 = loadCompleted_7 | _T_102202; // @[LoadQueue.scala 371:79:@44982.4]
  assign _T_102205 = allocatedEntries_8 == 1'h0; // @[LoadQueue.scala 371:82:@44983.4]
  assign _T_102206 = loadCompleted_8 | _T_102205; // @[LoadQueue.scala 371:79:@44984.4]
  assign _T_102208 = allocatedEntries_9 == 1'h0; // @[LoadQueue.scala 371:82:@44985.4]
  assign _T_102209 = loadCompleted_9 | _T_102208; // @[LoadQueue.scala 371:79:@44986.4]
  assign _T_102211 = allocatedEntries_10 == 1'h0; // @[LoadQueue.scala 371:82:@44987.4]
  assign _T_102212 = loadCompleted_10 | _T_102211; // @[LoadQueue.scala 371:79:@44988.4]
  assign _T_102214 = allocatedEntries_11 == 1'h0; // @[LoadQueue.scala 371:82:@44989.4]
  assign _T_102215 = loadCompleted_11 | _T_102214; // @[LoadQueue.scala 371:79:@44990.4]
  assign _T_102217 = allocatedEntries_12 == 1'h0; // @[LoadQueue.scala 371:82:@44991.4]
  assign _T_102218 = loadCompleted_12 | _T_102217; // @[LoadQueue.scala 371:79:@44992.4]
  assign _T_102220 = allocatedEntries_13 == 1'h0; // @[LoadQueue.scala 371:82:@44993.4]
  assign _T_102221 = loadCompleted_13 | _T_102220; // @[LoadQueue.scala 371:79:@44994.4]
  assign _T_102223 = allocatedEntries_14 == 1'h0; // @[LoadQueue.scala 371:82:@44995.4]
  assign _T_102224 = loadCompleted_14 | _T_102223; // @[LoadQueue.scala 371:79:@44996.4]
  assign _T_102226 = allocatedEntries_15 == 1'h0; // @[LoadQueue.scala 371:82:@44997.4]
  assign _T_102227 = loadCompleted_15 | _T_102226; // @[LoadQueue.scala 371:79:@44998.4]
  assign _T_102252 = _T_102182 & _T_102185; // @[LoadQueue.scala 371:96:@45017.4]
  assign _T_102253 = _T_102252 & _T_102188; // @[LoadQueue.scala 371:96:@45018.4]
  assign _T_102254 = _T_102253 & _T_102191; // @[LoadQueue.scala 371:96:@45019.4]
  assign _T_102255 = _T_102254 & _T_102194; // @[LoadQueue.scala 371:96:@45020.4]
  assign _T_102256 = _T_102255 & _T_102197; // @[LoadQueue.scala 371:96:@45021.4]
  assign _T_102257 = _T_102256 & _T_102200; // @[LoadQueue.scala 371:96:@45022.4]
  assign _T_102258 = _T_102257 & _T_102203; // @[LoadQueue.scala 371:96:@45023.4]
  assign _T_102259 = _T_102258 & _T_102206; // @[LoadQueue.scala 371:96:@45024.4]
  assign _T_102260 = _T_102259 & _T_102209; // @[LoadQueue.scala 371:96:@45025.4]
  assign _T_102261 = _T_102260 & _T_102212; // @[LoadQueue.scala 371:96:@45026.4]
  assign _T_102262 = _T_102261 & _T_102215; // @[LoadQueue.scala 371:96:@45027.4]
  assign _T_102263 = _T_102262 & _T_102218; // @[LoadQueue.scala 371:96:@45028.4]
  assign _T_102264 = _T_102263 & _T_102221; // @[LoadQueue.scala 371:96:@45029.4]
  assign _T_102265 = _T_102264 & _T_102224; // @[LoadQueue.scala 371:96:@45030.4]
  assign io_loadTail = tail; // @[LoadQueue.scala 380:15:@45034.4]
  assign io_loadHead = head; // @[LoadQueue.scala 379:15:@45033.4]
  assign io_loadEmpty = _T_102265 & _T_102227; // @[LoadQueue.scala 371:16:@45032.4]
  assign io_loadAddrDone_0 = addrKnown_0; // @[LoadQueue.scala 382:19:@45051.4]
  assign io_loadAddrDone_1 = addrKnown_1; // @[LoadQueue.scala 382:19:@45052.4]
  assign io_loadAddrDone_2 = addrKnown_2; // @[LoadQueue.scala 382:19:@45053.4]
  assign io_loadAddrDone_3 = addrKnown_3; // @[LoadQueue.scala 382:19:@45054.4]
  assign io_loadAddrDone_4 = addrKnown_4; // @[LoadQueue.scala 382:19:@45055.4]
  assign io_loadAddrDone_5 = addrKnown_5; // @[LoadQueue.scala 382:19:@45056.4]
  assign io_loadAddrDone_6 = addrKnown_6; // @[LoadQueue.scala 382:19:@45057.4]
  assign io_loadAddrDone_7 = addrKnown_7; // @[LoadQueue.scala 382:19:@45058.4]
  assign io_loadAddrDone_8 = addrKnown_8; // @[LoadQueue.scala 382:19:@45059.4]
  assign io_loadAddrDone_9 = addrKnown_9; // @[LoadQueue.scala 382:19:@45060.4]
  assign io_loadAddrDone_10 = addrKnown_10; // @[LoadQueue.scala 382:19:@45061.4]
  assign io_loadAddrDone_11 = addrKnown_11; // @[LoadQueue.scala 382:19:@45062.4]
  assign io_loadAddrDone_12 = addrKnown_12; // @[LoadQueue.scala 382:19:@45063.4]
  assign io_loadAddrDone_13 = addrKnown_13; // @[LoadQueue.scala 382:19:@45064.4]
  assign io_loadAddrDone_14 = addrKnown_14; // @[LoadQueue.scala 382:19:@45065.4]
  assign io_loadAddrDone_15 = addrKnown_15; // @[LoadQueue.scala 382:19:@45066.4]
  assign io_loadDataDone_0 = dataKnown_0; // @[LoadQueue.scala 383:19:@45067.4]
  assign io_loadDataDone_1 = dataKnown_1; // @[LoadQueue.scala 383:19:@45068.4]
  assign io_loadDataDone_2 = dataKnown_2; // @[LoadQueue.scala 383:19:@45069.4]
  assign io_loadDataDone_3 = dataKnown_3; // @[LoadQueue.scala 383:19:@45070.4]
  assign io_loadDataDone_4 = dataKnown_4; // @[LoadQueue.scala 383:19:@45071.4]
  assign io_loadDataDone_5 = dataKnown_5; // @[LoadQueue.scala 383:19:@45072.4]
  assign io_loadDataDone_6 = dataKnown_6; // @[LoadQueue.scala 383:19:@45073.4]
  assign io_loadDataDone_7 = dataKnown_7; // @[LoadQueue.scala 383:19:@45074.4]
  assign io_loadDataDone_8 = dataKnown_8; // @[LoadQueue.scala 383:19:@45075.4]
  assign io_loadDataDone_9 = dataKnown_9; // @[LoadQueue.scala 383:19:@45076.4]
  assign io_loadDataDone_10 = dataKnown_10; // @[LoadQueue.scala 383:19:@45077.4]
  assign io_loadDataDone_11 = dataKnown_11; // @[LoadQueue.scala 383:19:@45078.4]
  assign io_loadDataDone_12 = dataKnown_12; // @[LoadQueue.scala 383:19:@45079.4]
  assign io_loadDataDone_13 = dataKnown_13; // @[LoadQueue.scala 383:19:@45080.4]
  assign io_loadDataDone_14 = dataKnown_14; // @[LoadQueue.scala 383:19:@45081.4]
  assign io_loadDataDone_15 = dataKnown_15; // @[LoadQueue.scala 383:19:@45082.4]
  assign io_loadAddrQueue_0 = addrQ_0; // @[LoadQueue.scala 381:20:@45035.4]
  assign io_loadAddrQueue_1 = addrQ_1; // @[LoadQueue.scala 381:20:@45036.4]
  assign io_loadAddrQueue_2 = addrQ_2; // @[LoadQueue.scala 381:20:@45037.4]
  assign io_loadAddrQueue_3 = addrQ_3; // @[LoadQueue.scala 381:20:@45038.4]
  assign io_loadAddrQueue_4 = addrQ_4; // @[LoadQueue.scala 381:20:@45039.4]
  assign io_loadAddrQueue_5 = addrQ_5; // @[LoadQueue.scala 381:20:@45040.4]
  assign io_loadAddrQueue_6 = addrQ_6; // @[LoadQueue.scala 381:20:@45041.4]
  assign io_loadAddrQueue_7 = addrQ_7; // @[LoadQueue.scala 381:20:@45042.4]
  assign io_loadAddrQueue_8 = addrQ_8; // @[LoadQueue.scala 381:20:@45043.4]
  assign io_loadAddrQueue_9 = addrQ_9; // @[LoadQueue.scala 381:20:@45044.4]
  assign io_loadAddrQueue_10 = addrQ_10; // @[LoadQueue.scala 381:20:@45045.4]
  assign io_loadAddrQueue_11 = addrQ_11; // @[LoadQueue.scala 381:20:@45046.4]
  assign io_loadAddrQueue_12 = addrQ_12; // @[LoadQueue.scala 381:20:@45047.4]
  assign io_loadAddrQueue_13 = addrQ_13; // @[LoadQueue.scala 381:20:@45048.4]
  assign io_loadAddrQueue_14 = addrQ_14; // @[LoadQueue.scala 381:20:@45049.4]
  assign io_loadAddrQueue_15 = addrQ_15; // @[LoadQueue.scala 381:20:@45050.4]
  assign io_loadPorts_0_valid = _T_101984 | _T_101833; // @[LoadQueue.scala 350:38:@44842.6 LoadQueue.scala 353:38:@44846.6]
  assign io_loadPorts_0_bits = _T_101985 ? _GEN_2257 : 32'h0; // @[LoadQueue.scala 349:37:@44841.6 LoadQueue.scala 352:37:@44845.6]
  assign io_loadPorts_1_valid = _T_102124 | _T_101838; // @[LoadQueue.scala 350:38:@44946.6 LoadQueue.scala 353:38:@44950.6]
  assign io_loadPorts_1_bits = _T_102125 ? _GEN_2275 : 32'h0; // @[LoadQueue.scala 349:37:@44945.6 LoadQueue.scala 352:37:@44949.6]
  assign io_loadAddrToMem = _T_93618 ? _GEN_2047 : 32'h0; // @[LoadQueue.scala 248:24:@39139.6 LoadQueue.scala 251:24:@39143.6]
  assign io_loadEnableToMem = _T_93617 | loadRequest_15; // @[LoadQueue.scala 246:22:@39106.4 LoadQueue.scala 249:26:@39140.6 LoadQueue.scala 252:26:@39144.6]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  offsetQ_0 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  offsetQ_1 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  offsetQ_2 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  offsetQ_3 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  offsetQ_4 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  offsetQ_5 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  offsetQ_6 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  offsetQ_7 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  offsetQ_8 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  offsetQ_9 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  offsetQ_10 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  offsetQ_11 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  offsetQ_12 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  offsetQ_13 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  offsetQ_14 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  offsetQ_15 = _RAND_17[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  portQ_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  portQ_1 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  portQ_2 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  portQ_3 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  portQ_4 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  portQ_5 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  portQ_6 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  portQ_7 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  portQ_8 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  portQ_9 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  portQ_10 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  portQ_11 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  portQ_12 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  portQ_13 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  portQ_14 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  portQ_15 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  addrQ_0 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  addrQ_1 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  addrQ_2 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  addrQ_3 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  addrQ_4 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  addrQ_5 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  addrQ_6 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  addrQ_7 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  addrQ_8 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  addrQ_9 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  addrQ_10 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  addrQ_11 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  addrQ_12 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  addrQ_13 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  addrQ_14 = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  addrQ_15 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  dataQ_0 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  dataQ_1 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  dataQ_2 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  dataQ_3 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  dataQ_4 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  dataQ_5 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  dataQ_6 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  dataQ_7 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  dataQ_8 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  dataQ_9 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  dataQ_10 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  dataQ_11 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  dataQ_12 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  dataQ_13 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  dataQ_14 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  dataQ_15 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  addrKnown_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  addrKnown_1 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  addrKnown_2 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  addrKnown_3 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  addrKnown_4 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  addrKnown_5 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  addrKnown_6 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  addrKnown_7 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  addrKnown_8 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  addrKnown_9 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  addrKnown_10 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  addrKnown_11 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  addrKnown_12 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  addrKnown_13 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  addrKnown_14 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  addrKnown_15 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  dataKnown_0 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  dataKnown_1 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  dataKnown_2 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  dataKnown_3 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  dataKnown_4 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  dataKnown_5 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  dataKnown_6 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  dataKnown_7 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  dataKnown_8 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  dataKnown_9 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  dataKnown_10 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  dataKnown_11 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  dataKnown_12 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  dataKnown_13 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  dataKnown_14 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  dataKnown_15 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  loadCompleted_0 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  loadCompleted_1 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  loadCompleted_2 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  loadCompleted_3 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  loadCompleted_4 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  loadCompleted_5 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  loadCompleted_6 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  loadCompleted_7 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  loadCompleted_8 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  loadCompleted_9 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  loadCompleted_10 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  loadCompleted_11 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  loadCompleted_12 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  loadCompleted_13 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  loadCompleted_14 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  loadCompleted_15 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  allocatedEntries_0 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  allocatedEntries_1 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  allocatedEntries_2 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  allocatedEntries_3 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  allocatedEntries_4 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  allocatedEntries_5 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  allocatedEntries_6 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  allocatedEntries_7 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  allocatedEntries_8 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  allocatedEntries_9 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  allocatedEntries_10 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  allocatedEntries_11 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  allocatedEntries_12 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  allocatedEntries_13 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  allocatedEntries_14 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  allocatedEntries_15 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  bypassInitiated_0 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  bypassInitiated_1 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  bypassInitiated_2 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  bypassInitiated_3 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  bypassInitiated_4 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  bypassInitiated_5 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  bypassInitiated_6 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  bypassInitiated_7 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  bypassInitiated_8 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  bypassInitiated_9 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  bypassInitiated_10 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  bypassInitiated_11 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  bypassInitiated_12 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  bypassInitiated_13 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  bypassInitiated_14 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  bypassInitiated_15 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  checkBits_0 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  checkBits_1 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  checkBits_2 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  checkBits_3 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  checkBits_4 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  checkBits_5 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  checkBits_6 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  checkBits_7 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  checkBits_8 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  checkBits_9 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  checkBits_10 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  checkBits_11 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  checkBits_12 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  checkBits_13 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  checkBits_14 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  checkBits_15 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  previousStoreHead = _RAND_162[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  conflictPReg_0_0 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  conflictPReg_0_1 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  conflictPReg_0_2 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  conflictPReg_0_3 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  conflictPReg_0_4 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  conflictPReg_0_5 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  conflictPReg_0_6 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  conflictPReg_0_7 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  conflictPReg_0_8 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  conflictPReg_0_9 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  conflictPReg_0_10 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  conflictPReg_0_11 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  conflictPReg_0_12 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  conflictPReg_0_13 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  conflictPReg_0_14 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  conflictPReg_0_15 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  conflictPReg_1_0 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  conflictPReg_1_1 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  conflictPReg_1_2 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  conflictPReg_1_3 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  conflictPReg_1_4 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  conflictPReg_1_5 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  conflictPReg_1_6 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  conflictPReg_1_7 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  conflictPReg_1_8 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  conflictPReg_1_9 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  conflictPReg_1_10 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  conflictPReg_1_11 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  conflictPReg_1_12 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  conflictPReg_1_13 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  conflictPReg_1_14 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  conflictPReg_1_15 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  conflictPReg_2_0 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  conflictPReg_2_1 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  conflictPReg_2_2 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  conflictPReg_2_3 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  conflictPReg_2_4 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  conflictPReg_2_5 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  conflictPReg_2_6 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  conflictPReg_2_7 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  conflictPReg_2_8 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  conflictPReg_2_9 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  conflictPReg_2_10 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  conflictPReg_2_11 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  conflictPReg_2_12 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  conflictPReg_2_13 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  conflictPReg_2_14 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  conflictPReg_2_15 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  conflictPReg_3_0 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  conflictPReg_3_1 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  conflictPReg_3_2 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  conflictPReg_3_3 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  conflictPReg_3_4 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  conflictPReg_3_5 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  conflictPReg_3_6 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  conflictPReg_3_7 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  conflictPReg_3_8 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  conflictPReg_3_9 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  conflictPReg_3_10 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  conflictPReg_3_11 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  conflictPReg_3_12 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  conflictPReg_3_13 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  conflictPReg_3_14 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  conflictPReg_3_15 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  conflictPReg_4_0 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  conflictPReg_4_1 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  conflictPReg_4_2 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  conflictPReg_4_3 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  conflictPReg_4_4 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  conflictPReg_4_5 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  conflictPReg_4_6 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  conflictPReg_4_7 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  conflictPReg_4_8 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  conflictPReg_4_9 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  conflictPReg_4_10 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  conflictPReg_4_11 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  conflictPReg_4_12 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  conflictPReg_4_13 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  conflictPReg_4_14 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  conflictPReg_4_15 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  conflictPReg_5_0 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  conflictPReg_5_1 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  conflictPReg_5_2 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  conflictPReg_5_3 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  conflictPReg_5_4 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  conflictPReg_5_5 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  conflictPReg_5_6 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  conflictPReg_5_7 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  conflictPReg_5_8 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  conflictPReg_5_9 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  conflictPReg_5_10 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  conflictPReg_5_11 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  conflictPReg_5_12 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  conflictPReg_5_13 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  conflictPReg_5_14 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  conflictPReg_5_15 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  conflictPReg_6_0 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  conflictPReg_6_1 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  conflictPReg_6_2 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  conflictPReg_6_3 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  conflictPReg_6_4 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  conflictPReg_6_5 = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  conflictPReg_6_6 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  conflictPReg_6_7 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  conflictPReg_6_8 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  conflictPReg_6_9 = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  conflictPReg_6_10 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  conflictPReg_6_11 = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  conflictPReg_6_12 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  conflictPReg_6_13 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  conflictPReg_6_14 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  conflictPReg_6_15 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  conflictPReg_7_0 = _RAND_275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  conflictPReg_7_1 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  conflictPReg_7_2 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  conflictPReg_7_3 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  conflictPReg_7_4 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  conflictPReg_7_5 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  conflictPReg_7_6 = _RAND_281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  conflictPReg_7_7 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  conflictPReg_7_8 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  conflictPReg_7_9 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  conflictPReg_7_10 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  conflictPReg_7_11 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  conflictPReg_7_12 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  conflictPReg_7_13 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  conflictPReg_7_14 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  conflictPReg_7_15 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  conflictPReg_8_0 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  conflictPReg_8_1 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  conflictPReg_8_2 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  conflictPReg_8_3 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  conflictPReg_8_4 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  conflictPReg_8_5 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  conflictPReg_8_6 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  conflictPReg_8_7 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  conflictPReg_8_8 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  conflictPReg_8_9 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  conflictPReg_8_10 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  conflictPReg_8_11 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  conflictPReg_8_12 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  conflictPReg_8_13 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  conflictPReg_8_14 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  conflictPReg_8_15 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  conflictPReg_9_0 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  conflictPReg_9_1 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  conflictPReg_9_2 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  conflictPReg_9_3 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  conflictPReg_9_4 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  conflictPReg_9_5 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  conflictPReg_9_6 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  conflictPReg_9_7 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  conflictPReg_9_8 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  conflictPReg_9_9 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  conflictPReg_9_10 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  conflictPReg_9_11 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  conflictPReg_9_12 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  conflictPReg_9_13 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  conflictPReg_9_14 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  conflictPReg_9_15 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  conflictPReg_10_0 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  conflictPReg_10_1 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  conflictPReg_10_2 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  conflictPReg_10_3 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  conflictPReg_10_4 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  conflictPReg_10_5 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  conflictPReg_10_6 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  conflictPReg_10_7 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  conflictPReg_10_8 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  conflictPReg_10_9 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  conflictPReg_10_10 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  conflictPReg_10_11 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  conflictPReg_10_12 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  conflictPReg_10_13 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  conflictPReg_10_14 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  conflictPReg_10_15 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  conflictPReg_11_0 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  conflictPReg_11_1 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  conflictPReg_11_2 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  conflictPReg_11_3 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  conflictPReg_11_4 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  conflictPReg_11_5 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  conflictPReg_11_6 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  conflictPReg_11_7 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  conflictPReg_11_8 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  conflictPReg_11_9 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  conflictPReg_11_10 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  conflictPReg_11_11 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  conflictPReg_11_12 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  conflictPReg_11_13 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  conflictPReg_11_14 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  conflictPReg_11_15 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  conflictPReg_12_0 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  conflictPReg_12_1 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  conflictPReg_12_2 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  conflictPReg_12_3 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  conflictPReg_12_4 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  conflictPReg_12_5 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  conflictPReg_12_6 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  conflictPReg_12_7 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  conflictPReg_12_8 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  conflictPReg_12_9 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  conflictPReg_12_10 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  conflictPReg_12_11 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  conflictPReg_12_12 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  conflictPReg_12_13 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  conflictPReg_12_14 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  conflictPReg_12_15 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  conflictPReg_13_0 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  conflictPReg_13_1 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  conflictPReg_13_2 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  conflictPReg_13_3 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  conflictPReg_13_4 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  conflictPReg_13_5 = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  conflictPReg_13_6 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  conflictPReg_13_7 = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  conflictPReg_13_8 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  conflictPReg_13_9 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  conflictPReg_13_10 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  conflictPReg_13_11 = _RAND_382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  conflictPReg_13_12 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  conflictPReg_13_13 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  conflictPReg_13_14 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  conflictPReg_13_15 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  conflictPReg_14_0 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  conflictPReg_14_1 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  conflictPReg_14_2 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  conflictPReg_14_3 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  conflictPReg_14_4 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  conflictPReg_14_5 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  conflictPReg_14_6 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  conflictPReg_14_7 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  conflictPReg_14_8 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  conflictPReg_14_9 = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  conflictPReg_14_10 = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  conflictPReg_14_11 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  conflictPReg_14_12 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  conflictPReg_14_13 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  conflictPReg_14_14 = _RAND_401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  conflictPReg_14_15 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  conflictPReg_15_0 = _RAND_403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  conflictPReg_15_1 = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  conflictPReg_15_2 = _RAND_405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  conflictPReg_15_3 = _RAND_406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  conflictPReg_15_4 = _RAND_407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  conflictPReg_15_5 = _RAND_408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  conflictPReg_15_6 = _RAND_409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  conflictPReg_15_7 = _RAND_410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  conflictPReg_15_8 = _RAND_411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  conflictPReg_15_9 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  conflictPReg_15_10 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  conflictPReg_15_11 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  conflictPReg_15_12 = _RAND_415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  conflictPReg_15_13 = _RAND_416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  conflictPReg_15_14 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  conflictPReg_15_15 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_0 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_1 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_2 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_3 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_4 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_5 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_6 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_7 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_8 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_9 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_10 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_11 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_12 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_13 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_14 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_15 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_0 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_1 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_2 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_3 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_4 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_5 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_6 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_7 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_8 = _RAND_443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_9 = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_10 = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_11 = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_12 = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_13 = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_14 = _RAND_449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_15 = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_0 = _RAND_451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_1 = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_2 = _RAND_453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_3 = _RAND_454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_4 = _RAND_455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_5 = _RAND_456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_6 = _RAND_457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_7 = _RAND_458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_8 = _RAND_459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_9 = _RAND_460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_10 = _RAND_461[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_11 = _RAND_462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_12 = _RAND_463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_13 = _RAND_464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_14 = _RAND_465[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_15 = _RAND_466[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_0 = _RAND_467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_1 = _RAND_468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_2 = _RAND_469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_3 = _RAND_470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_4 = _RAND_471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_5 = _RAND_472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_6 = _RAND_473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_7 = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_8 = _RAND_475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_9 = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_10 = _RAND_477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_11 = _RAND_478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_12 = _RAND_479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_13 = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_14 = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_15 = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_0 = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_1 = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_2 = _RAND_485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_3 = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_4 = _RAND_487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_5 = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_6 = _RAND_489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_7 = _RAND_490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_8 = _RAND_491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_9 = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_10 = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_11 = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_12 = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_13 = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_14 = _RAND_497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_15 = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_0 = _RAND_499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_1 = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_2 = _RAND_501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_3 = _RAND_502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_4 = _RAND_503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_5 = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_6 = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_7 = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_8 = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_9 = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_10 = _RAND_509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_11 = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_12 = _RAND_511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_13 = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_14 = _RAND_513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_15 = _RAND_514[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_0 = _RAND_515[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_1 = _RAND_516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_2 = _RAND_517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_3 = _RAND_518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_4 = _RAND_519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_5 = _RAND_520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_6 = _RAND_521[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_7 = _RAND_522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_8 = _RAND_523[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_9 = _RAND_524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_10 = _RAND_525[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_11 = _RAND_526[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_12 = _RAND_527[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_13 = _RAND_528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_14 = _RAND_529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_15 = _RAND_530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_0 = _RAND_531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_1 = _RAND_532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_2 = _RAND_533[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_3 = _RAND_534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_4 = _RAND_535[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_5 = _RAND_536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_6 = _RAND_537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_7 = _RAND_538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_8 = _RAND_539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_9 = _RAND_540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_10 = _RAND_541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_11 = _RAND_542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_12 = _RAND_543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_13 = _RAND_544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_14 = _RAND_545[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_15 = _RAND_546[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_0 = _RAND_547[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_1 = _RAND_548[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_2 = _RAND_549[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_3 = _RAND_550[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_4 = _RAND_551[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_5 = _RAND_552[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_6 = _RAND_553[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_7 = _RAND_554[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_8 = _RAND_555[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_9 = _RAND_556[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_10 = _RAND_557[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_11 = _RAND_558[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_12 = _RAND_559[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_13 = _RAND_560[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_14 = _RAND_561[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_15 = _RAND_562[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_0 = _RAND_563[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_1 = _RAND_564[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_2 = _RAND_565[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_3 = _RAND_566[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_4 = _RAND_567[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_5 = _RAND_568[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_6 = _RAND_569[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_7 = _RAND_570[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_8 = _RAND_571[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_9 = _RAND_572[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_10 = _RAND_573[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_11 = _RAND_574[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_12 = _RAND_575[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_13 = _RAND_576[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_14 = _RAND_577[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_15 = _RAND_578[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_0 = _RAND_579[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_1 = _RAND_580[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_2 = _RAND_581[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_3 = _RAND_582[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_4 = _RAND_583[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_5 = _RAND_584[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_6 = _RAND_585[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_7 = _RAND_586[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_8 = _RAND_587[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_9 = _RAND_588[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_10 = _RAND_589[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_11 = _RAND_590[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_12 = _RAND_591[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_13 = _RAND_592[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_14 = _RAND_593[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_15 = _RAND_594[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_0 = _RAND_595[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_1 = _RAND_596[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_2 = _RAND_597[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_3 = _RAND_598[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_4 = _RAND_599[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_5 = _RAND_600[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_6 = _RAND_601[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_7 = _RAND_602[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_8 = _RAND_603[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_9 = _RAND_604[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_10 = _RAND_605[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_11 = _RAND_606[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_12 = _RAND_607[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_13 = _RAND_608[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_14 = _RAND_609[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_15 = _RAND_610[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_0 = _RAND_611[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_1 = _RAND_612[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_2 = _RAND_613[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_3 = _RAND_614[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_4 = _RAND_615[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_5 = _RAND_616[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_6 = _RAND_617[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_7 = _RAND_618[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_8 = _RAND_619[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_9 = _RAND_620[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_10 = _RAND_621[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_11 = _RAND_622[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_12 = _RAND_623[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_13 = _RAND_624[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_14 = _RAND_625[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_15 = _RAND_626[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_0 = _RAND_627[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_1 = _RAND_628[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_2 = _RAND_629[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_3 = _RAND_630[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_4 = _RAND_631[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_5 = _RAND_632[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_6 = _RAND_633[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_7 = _RAND_634[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_8 = _RAND_635[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_9 = _RAND_636[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_10 = _RAND_637[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_11 = _RAND_638[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_12 = _RAND_639[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_13 = _RAND_640[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_14 = _RAND_641[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_15 = _RAND_642[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_0 = _RAND_643[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_1 = _RAND_644[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_2 = _RAND_645[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_3 = _RAND_646[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_4 = _RAND_647[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_5 = _RAND_648[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_6 = _RAND_649[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_7 = _RAND_650[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_8 = _RAND_651[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_9 = _RAND_652[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_10 = _RAND_653[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_11 = _RAND_654[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_12 = _RAND_655[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_13 = _RAND_656[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_14 = _RAND_657[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_15 = _RAND_658[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_0 = _RAND_659[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_1 = _RAND_660[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_2 = _RAND_661[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_3 = _RAND_662[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_4 = _RAND_663[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_5 = _RAND_664[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_6 = _RAND_665[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_7 = _RAND_666[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_8 = _RAND_667[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_9 = _RAND_668[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_10 = _RAND_669[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_11 = _RAND_670[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_12 = _RAND_671[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_13 = _RAND_672[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_14 = _RAND_673[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_15 = _RAND_674[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_0 = _RAND_675[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_1 = _RAND_676[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_2 = _RAND_677[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_3 = _RAND_678[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_4 = _RAND_679[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_5 = _RAND_680[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_6 = _RAND_681[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_7 = _RAND_682[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_8 = _RAND_683[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_9 = _RAND_684[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_10 = _RAND_685[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_11 = _RAND_686[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_12 = _RAND_687[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_13 = _RAND_688[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_14 = _RAND_689[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_15 = _RAND_690[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{`RANDOM}};
  shiftedStoreDataQPreg_0 = _RAND_691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{`RANDOM}};
  shiftedStoreDataQPreg_1 = _RAND_692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{`RANDOM}};
  shiftedStoreDataQPreg_2 = _RAND_693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{`RANDOM}};
  shiftedStoreDataQPreg_3 = _RAND_694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{`RANDOM}};
  shiftedStoreDataQPreg_4 = _RAND_695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{`RANDOM}};
  shiftedStoreDataQPreg_5 = _RAND_696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{`RANDOM}};
  shiftedStoreDataQPreg_6 = _RAND_697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{`RANDOM}};
  shiftedStoreDataQPreg_7 = _RAND_698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{`RANDOM}};
  shiftedStoreDataQPreg_8 = _RAND_699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{`RANDOM}};
  shiftedStoreDataQPreg_9 = _RAND_700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{`RANDOM}};
  shiftedStoreDataQPreg_10 = _RAND_701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{`RANDOM}};
  shiftedStoreDataQPreg_11 = _RAND_702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{`RANDOM}};
  shiftedStoreDataQPreg_12 = _RAND_703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{`RANDOM}};
  shiftedStoreDataQPreg_13 = _RAND_704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{`RANDOM}};
  shiftedStoreDataQPreg_14 = _RAND_705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{`RANDOM}};
  shiftedStoreDataQPreg_15 = _RAND_706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{`RANDOM}};
  addrKnownPReg_0 = _RAND_707[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{`RANDOM}};
  addrKnownPReg_1 = _RAND_708[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{`RANDOM}};
  addrKnownPReg_2 = _RAND_709[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{`RANDOM}};
  addrKnownPReg_3 = _RAND_710[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{`RANDOM}};
  addrKnownPReg_4 = _RAND_711[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{`RANDOM}};
  addrKnownPReg_5 = _RAND_712[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{`RANDOM}};
  addrKnownPReg_6 = _RAND_713[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{`RANDOM}};
  addrKnownPReg_7 = _RAND_714[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{`RANDOM}};
  addrKnownPReg_8 = _RAND_715[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{`RANDOM}};
  addrKnownPReg_9 = _RAND_716[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{`RANDOM}};
  addrKnownPReg_10 = _RAND_717[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{`RANDOM}};
  addrKnownPReg_11 = _RAND_718[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{`RANDOM}};
  addrKnownPReg_12 = _RAND_719[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{`RANDOM}};
  addrKnownPReg_13 = _RAND_720[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{`RANDOM}};
  addrKnownPReg_14 = _RAND_721[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{`RANDOM}};
  addrKnownPReg_15 = _RAND_722[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{`RANDOM}};
  dataKnownPReg_0 = _RAND_723[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{`RANDOM}};
  dataKnownPReg_1 = _RAND_724[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{`RANDOM}};
  dataKnownPReg_2 = _RAND_725[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{`RANDOM}};
  dataKnownPReg_3 = _RAND_726[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{`RANDOM}};
  dataKnownPReg_4 = _RAND_727[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{`RANDOM}};
  dataKnownPReg_5 = _RAND_728[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{`RANDOM}};
  dataKnownPReg_6 = _RAND_729[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{`RANDOM}};
  dataKnownPReg_7 = _RAND_730[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{`RANDOM}};
  dataKnownPReg_8 = _RAND_731[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{`RANDOM}};
  dataKnownPReg_9 = _RAND_732[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{`RANDOM}};
  dataKnownPReg_10 = _RAND_733[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{`RANDOM}};
  dataKnownPReg_11 = _RAND_734[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{`RANDOM}};
  dataKnownPReg_12 = _RAND_735[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{`RANDOM}};
  dataKnownPReg_13 = _RAND_736[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{`RANDOM}};
  dataKnownPReg_14 = _RAND_737[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{`RANDOM}};
  dataKnownPReg_15 = _RAND_738[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{`RANDOM}};
  prevPriorityRequest_15 = _RAND_739[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{`RANDOM}};
  prevPriorityRequest_14 = _RAND_740[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{`RANDOM}};
  prevPriorityRequest_13 = _RAND_741[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{`RANDOM}};
  prevPriorityRequest_12 = _RAND_742[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{`RANDOM}};
  prevPriorityRequest_11 = _RAND_743[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{`RANDOM}};
  prevPriorityRequest_10 = _RAND_744[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{`RANDOM}};
  prevPriorityRequest_9 = _RAND_745[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{`RANDOM}};
  prevPriorityRequest_8 = _RAND_746[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{`RANDOM}};
  prevPriorityRequest_7 = _RAND_747[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{`RANDOM}};
  prevPriorityRequest_6 = _RAND_748[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{`RANDOM}};
  prevPriorityRequest_5 = _RAND_749[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{`RANDOM}};
  prevPriorityRequest_4 = _RAND_750[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{`RANDOM}};
  prevPriorityRequest_3 = _RAND_751[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{`RANDOM}};
  prevPriorityRequest_2 = _RAND_752[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_753 = {1{`RANDOM}};
  prevPriorityRequest_1 = _RAND_753[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_754 = {1{`RANDOM}};
  prevPriorityRequest_0 = _RAND_754[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      head <= 4'h0;
    end else begin
      head <= _GEN_2310[3:0];
    end
    if (reset) begin
      tail <= 4'h0;
    end else begin
      tail <= _GEN_2311[3:0];
    end
    if (reset) begin
      offsetQ_0 <= 4'h0;
    end else begin
      if (initBits_0) begin
        if (4'hf == _T_1932) begin
          offsetQ_0 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1932) begin
            offsetQ_0 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1932) begin
              offsetQ_0 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1932) begin
                offsetQ_0 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1932) begin
                  offsetQ_0 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1932) begin
                    offsetQ_0 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1932) begin
                      offsetQ_0 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1932) begin
                        offsetQ_0 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1932) begin
                          offsetQ_0 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1932) begin
                            offsetQ_0 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1932) begin
                              offsetQ_0 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1932) begin
                                offsetQ_0 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1932) begin
                                  offsetQ_0 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1932) begin
                                    offsetQ_0 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1932) begin
                                      offsetQ_0 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_0 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_1 <= 4'h0;
    end else begin
      if (initBits_1) begin
        if (4'hf == _T_1950) begin
          offsetQ_1 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1950) begin
            offsetQ_1 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1950) begin
              offsetQ_1 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1950) begin
                offsetQ_1 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1950) begin
                  offsetQ_1 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1950) begin
                    offsetQ_1 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1950) begin
                      offsetQ_1 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1950) begin
                        offsetQ_1 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1950) begin
                          offsetQ_1 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1950) begin
                            offsetQ_1 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1950) begin
                              offsetQ_1 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1950) begin
                                offsetQ_1 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1950) begin
                                  offsetQ_1 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1950) begin
                                    offsetQ_1 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1950) begin
                                      offsetQ_1 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_1 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_2 <= 4'h0;
    end else begin
      if (initBits_2) begin
        if (4'hf == _T_1968) begin
          offsetQ_2 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1968) begin
            offsetQ_2 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1968) begin
              offsetQ_2 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1968) begin
                offsetQ_2 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1968) begin
                  offsetQ_2 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1968) begin
                    offsetQ_2 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1968) begin
                      offsetQ_2 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1968) begin
                        offsetQ_2 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1968) begin
                          offsetQ_2 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1968) begin
                            offsetQ_2 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1968) begin
                              offsetQ_2 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1968) begin
                                offsetQ_2 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1968) begin
                                  offsetQ_2 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1968) begin
                                    offsetQ_2 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1968) begin
                                      offsetQ_2 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_2 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_3 <= 4'h0;
    end else begin
      if (initBits_3) begin
        if (4'hf == _T_1986) begin
          offsetQ_3 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1986) begin
            offsetQ_3 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1986) begin
              offsetQ_3 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1986) begin
                offsetQ_3 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1986) begin
                  offsetQ_3 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1986) begin
                    offsetQ_3 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1986) begin
                      offsetQ_3 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1986) begin
                        offsetQ_3 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1986) begin
                          offsetQ_3 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1986) begin
                            offsetQ_3 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1986) begin
                              offsetQ_3 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1986) begin
                                offsetQ_3 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1986) begin
                                  offsetQ_3 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1986) begin
                                    offsetQ_3 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1986) begin
                                      offsetQ_3 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_3 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_4 <= 4'h0;
    end else begin
      if (initBits_4) begin
        if (4'hf == _T_2004) begin
          offsetQ_4 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2004) begin
            offsetQ_4 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2004) begin
              offsetQ_4 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2004) begin
                offsetQ_4 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2004) begin
                  offsetQ_4 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2004) begin
                    offsetQ_4 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2004) begin
                      offsetQ_4 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2004) begin
                        offsetQ_4 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2004) begin
                          offsetQ_4 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2004) begin
                            offsetQ_4 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2004) begin
                              offsetQ_4 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2004) begin
                                offsetQ_4 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2004) begin
                                  offsetQ_4 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2004) begin
                                    offsetQ_4 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2004) begin
                                      offsetQ_4 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_4 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_5 <= 4'h0;
    end else begin
      if (initBits_5) begin
        if (4'hf == _T_2022) begin
          offsetQ_5 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2022) begin
            offsetQ_5 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2022) begin
              offsetQ_5 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2022) begin
                offsetQ_5 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2022) begin
                  offsetQ_5 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2022) begin
                    offsetQ_5 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2022) begin
                      offsetQ_5 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2022) begin
                        offsetQ_5 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2022) begin
                          offsetQ_5 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2022) begin
                            offsetQ_5 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2022) begin
                              offsetQ_5 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2022) begin
                                offsetQ_5 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2022) begin
                                  offsetQ_5 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2022) begin
                                    offsetQ_5 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2022) begin
                                      offsetQ_5 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_5 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_6 <= 4'h0;
    end else begin
      if (initBits_6) begin
        if (4'hf == _T_2040) begin
          offsetQ_6 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2040) begin
            offsetQ_6 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2040) begin
              offsetQ_6 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2040) begin
                offsetQ_6 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2040) begin
                  offsetQ_6 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2040) begin
                    offsetQ_6 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2040) begin
                      offsetQ_6 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2040) begin
                        offsetQ_6 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2040) begin
                          offsetQ_6 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2040) begin
                            offsetQ_6 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2040) begin
                              offsetQ_6 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2040) begin
                                offsetQ_6 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2040) begin
                                  offsetQ_6 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2040) begin
                                    offsetQ_6 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2040) begin
                                      offsetQ_6 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_6 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_7 <= 4'h0;
    end else begin
      if (initBits_7) begin
        if (4'hf == _T_2058) begin
          offsetQ_7 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2058) begin
            offsetQ_7 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2058) begin
              offsetQ_7 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2058) begin
                offsetQ_7 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2058) begin
                  offsetQ_7 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2058) begin
                    offsetQ_7 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2058) begin
                      offsetQ_7 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2058) begin
                        offsetQ_7 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2058) begin
                          offsetQ_7 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2058) begin
                            offsetQ_7 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2058) begin
                              offsetQ_7 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2058) begin
                                offsetQ_7 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2058) begin
                                  offsetQ_7 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2058) begin
                                    offsetQ_7 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2058) begin
                                      offsetQ_7 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_7 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_8 <= 4'h0;
    end else begin
      if (initBits_8) begin
        if (4'hf == _T_2076) begin
          offsetQ_8 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2076) begin
            offsetQ_8 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2076) begin
              offsetQ_8 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2076) begin
                offsetQ_8 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2076) begin
                  offsetQ_8 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2076) begin
                    offsetQ_8 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2076) begin
                      offsetQ_8 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2076) begin
                        offsetQ_8 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2076) begin
                          offsetQ_8 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2076) begin
                            offsetQ_8 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2076) begin
                              offsetQ_8 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2076) begin
                                offsetQ_8 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2076) begin
                                  offsetQ_8 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2076) begin
                                    offsetQ_8 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2076) begin
                                      offsetQ_8 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_8 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_9 <= 4'h0;
    end else begin
      if (initBits_9) begin
        if (4'hf == _T_2094) begin
          offsetQ_9 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2094) begin
            offsetQ_9 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2094) begin
              offsetQ_9 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2094) begin
                offsetQ_9 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2094) begin
                  offsetQ_9 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2094) begin
                    offsetQ_9 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2094) begin
                      offsetQ_9 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2094) begin
                        offsetQ_9 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2094) begin
                          offsetQ_9 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2094) begin
                            offsetQ_9 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2094) begin
                              offsetQ_9 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2094) begin
                                offsetQ_9 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2094) begin
                                  offsetQ_9 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2094) begin
                                    offsetQ_9 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2094) begin
                                      offsetQ_9 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_9 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_10 <= 4'h0;
    end else begin
      if (initBits_10) begin
        if (4'hf == _T_2112) begin
          offsetQ_10 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2112) begin
            offsetQ_10 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2112) begin
              offsetQ_10 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2112) begin
                offsetQ_10 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2112) begin
                  offsetQ_10 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2112) begin
                    offsetQ_10 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2112) begin
                      offsetQ_10 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2112) begin
                        offsetQ_10 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2112) begin
                          offsetQ_10 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2112) begin
                            offsetQ_10 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2112) begin
                              offsetQ_10 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2112) begin
                                offsetQ_10 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2112) begin
                                  offsetQ_10 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2112) begin
                                    offsetQ_10 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2112) begin
                                      offsetQ_10 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_10 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_11 <= 4'h0;
    end else begin
      if (initBits_11) begin
        if (4'hf == _T_2130) begin
          offsetQ_11 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2130) begin
            offsetQ_11 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2130) begin
              offsetQ_11 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2130) begin
                offsetQ_11 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2130) begin
                  offsetQ_11 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2130) begin
                    offsetQ_11 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2130) begin
                      offsetQ_11 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2130) begin
                        offsetQ_11 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2130) begin
                          offsetQ_11 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2130) begin
                            offsetQ_11 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2130) begin
                              offsetQ_11 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2130) begin
                                offsetQ_11 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2130) begin
                                  offsetQ_11 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2130) begin
                                    offsetQ_11 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2130) begin
                                      offsetQ_11 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_11 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_12 <= 4'h0;
    end else begin
      if (initBits_12) begin
        if (4'hf == _T_2148) begin
          offsetQ_12 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2148) begin
            offsetQ_12 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2148) begin
              offsetQ_12 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2148) begin
                offsetQ_12 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2148) begin
                  offsetQ_12 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2148) begin
                    offsetQ_12 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2148) begin
                      offsetQ_12 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2148) begin
                        offsetQ_12 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2148) begin
                          offsetQ_12 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2148) begin
                            offsetQ_12 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2148) begin
                              offsetQ_12 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2148) begin
                                offsetQ_12 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2148) begin
                                  offsetQ_12 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2148) begin
                                    offsetQ_12 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2148) begin
                                      offsetQ_12 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_12 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_13 <= 4'h0;
    end else begin
      if (initBits_13) begin
        if (4'hf == _T_2166) begin
          offsetQ_13 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2166) begin
            offsetQ_13 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2166) begin
              offsetQ_13 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2166) begin
                offsetQ_13 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2166) begin
                  offsetQ_13 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2166) begin
                    offsetQ_13 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2166) begin
                      offsetQ_13 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2166) begin
                        offsetQ_13 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2166) begin
                          offsetQ_13 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2166) begin
                            offsetQ_13 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2166) begin
                              offsetQ_13 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2166) begin
                                offsetQ_13 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2166) begin
                                  offsetQ_13 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2166) begin
                                    offsetQ_13 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2166) begin
                                      offsetQ_13 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_13 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_14 <= 4'h0;
    end else begin
      if (initBits_14) begin
        if (4'hf == _T_2184) begin
          offsetQ_14 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2184) begin
            offsetQ_14 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2184) begin
              offsetQ_14 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2184) begin
                offsetQ_14 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2184) begin
                  offsetQ_14 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2184) begin
                    offsetQ_14 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2184) begin
                      offsetQ_14 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2184) begin
                        offsetQ_14 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2184) begin
                          offsetQ_14 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2184) begin
                            offsetQ_14 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2184) begin
                              offsetQ_14 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2184) begin
                                offsetQ_14 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2184) begin
                                  offsetQ_14 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2184) begin
                                    offsetQ_14 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2184) begin
                                      offsetQ_14 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_14 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_15 <= 4'h0;
    end else begin
      if (initBits_15) begin
        if (4'hf == _T_2202) begin
          offsetQ_15 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2202) begin
            offsetQ_15 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2202) begin
              offsetQ_15 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2202) begin
                offsetQ_15 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2202) begin
                  offsetQ_15 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2202) begin
                    offsetQ_15 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2202) begin
                      offsetQ_15 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2202) begin
                        offsetQ_15 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2202) begin
                          offsetQ_15 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2202) begin
                            offsetQ_15 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2202) begin
                              offsetQ_15 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2202) begin
                                offsetQ_15 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2202) begin
                                  offsetQ_15 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2202) begin
                                    offsetQ_15 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2202) begin
                                      offsetQ_15 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_15 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        if (4'hf == _T_1932) begin
          portQ_0 <= 1'h0;
        end else begin
          if (4'he == _T_1932) begin
            portQ_0 <= 1'h0;
          end else begin
            if (4'hd == _T_1932) begin
              portQ_0 <= 1'h0;
            end else begin
              if (4'hc == _T_1932) begin
                portQ_0 <= 1'h0;
              end else begin
                if (4'hb == _T_1932) begin
                  portQ_0 <= 1'h0;
                end else begin
                  if (4'ha == _T_1932) begin
                    portQ_0 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_1932) begin
                      portQ_0 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_1932) begin
                        portQ_0 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_1932) begin
                          portQ_0 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_1932) begin
                            portQ_0 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_1932) begin
                              portQ_0 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_1932) begin
                                portQ_0 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_1932) begin
                                  portQ_0 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_1932) begin
                                    portQ_0 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_1932) begin
                                      portQ_0 <= io_bbLoadPorts_1;
                                    end else begin
                                      portQ_0 <= 1'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        if (4'hf == _T_1950) begin
          portQ_1 <= 1'h0;
        end else begin
          if (4'he == _T_1950) begin
            portQ_1 <= 1'h0;
          end else begin
            if (4'hd == _T_1950) begin
              portQ_1 <= 1'h0;
            end else begin
              if (4'hc == _T_1950) begin
                portQ_1 <= 1'h0;
              end else begin
                if (4'hb == _T_1950) begin
                  portQ_1 <= 1'h0;
                end else begin
                  if (4'ha == _T_1950) begin
                    portQ_1 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_1950) begin
                      portQ_1 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_1950) begin
                        portQ_1 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_1950) begin
                          portQ_1 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_1950) begin
                            portQ_1 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_1950) begin
                              portQ_1 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_1950) begin
                                portQ_1 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_1950) begin
                                  portQ_1 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_1950) begin
                                    portQ_1 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_1950) begin
                                      portQ_1 <= io_bbLoadPorts_1;
                                    end else begin
                                      portQ_1 <= 1'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        if (4'hf == _T_1968) begin
          portQ_2 <= 1'h0;
        end else begin
          if (4'he == _T_1968) begin
            portQ_2 <= 1'h0;
          end else begin
            if (4'hd == _T_1968) begin
              portQ_2 <= 1'h0;
            end else begin
              if (4'hc == _T_1968) begin
                portQ_2 <= 1'h0;
              end else begin
                if (4'hb == _T_1968) begin
                  portQ_2 <= 1'h0;
                end else begin
                  if (4'ha == _T_1968) begin
                    portQ_2 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_1968) begin
                      portQ_2 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_1968) begin
                        portQ_2 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_1968) begin
                          portQ_2 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_1968) begin
                            portQ_2 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_1968) begin
                              portQ_2 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_1968) begin
                                portQ_2 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_1968) begin
                                  portQ_2 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_1968) begin
                                    portQ_2 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_1968) begin
                                      portQ_2 <= io_bbLoadPorts_1;
                                    end else begin
                                      portQ_2 <= 1'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        if (4'hf == _T_1986) begin
          portQ_3 <= 1'h0;
        end else begin
          if (4'he == _T_1986) begin
            portQ_3 <= 1'h0;
          end else begin
            if (4'hd == _T_1986) begin
              portQ_3 <= 1'h0;
            end else begin
              if (4'hc == _T_1986) begin
                portQ_3 <= 1'h0;
              end else begin
                if (4'hb == _T_1986) begin
                  portQ_3 <= 1'h0;
                end else begin
                  if (4'ha == _T_1986) begin
                    portQ_3 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_1986) begin
                      portQ_3 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_1986) begin
                        portQ_3 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_1986) begin
                          portQ_3 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_1986) begin
                            portQ_3 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_1986) begin
                              portQ_3 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_1986) begin
                                portQ_3 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_1986) begin
                                  portQ_3 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_1986) begin
                                    portQ_3 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_1986) begin
                                      portQ_3 <= io_bbLoadPorts_1;
                                    end else begin
                                      portQ_3 <= 1'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        if (4'hf == _T_2004) begin
          portQ_4 <= 1'h0;
        end else begin
          if (4'he == _T_2004) begin
            portQ_4 <= 1'h0;
          end else begin
            if (4'hd == _T_2004) begin
              portQ_4 <= 1'h0;
            end else begin
              if (4'hc == _T_2004) begin
                portQ_4 <= 1'h0;
              end else begin
                if (4'hb == _T_2004) begin
                  portQ_4 <= 1'h0;
                end else begin
                  if (4'ha == _T_2004) begin
                    portQ_4 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_2004) begin
                      portQ_4 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_2004) begin
                        portQ_4 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_2004) begin
                          portQ_4 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_2004) begin
                            portQ_4 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_2004) begin
                              portQ_4 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_2004) begin
                                portQ_4 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_2004) begin
                                  portQ_4 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_2004) begin
                                    portQ_4 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_2004) begin
                                      portQ_4 <= io_bbLoadPorts_1;
                                    end else begin
                                      portQ_4 <= 1'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        if (4'hf == _T_2022) begin
          portQ_5 <= 1'h0;
        end else begin
          if (4'he == _T_2022) begin
            portQ_5 <= 1'h0;
          end else begin
            if (4'hd == _T_2022) begin
              portQ_5 <= 1'h0;
            end else begin
              if (4'hc == _T_2022) begin
                portQ_5 <= 1'h0;
              end else begin
                if (4'hb == _T_2022) begin
                  portQ_5 <= 1'h0;
                end else begin
                  if (4'ha == _T_2022) begin
                    portQ_5 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_2022) begin
                      portQ_5 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_2022) begin
                        portQ_5 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_2022) begin
                          portQ_5 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_2022) begin
                            portQ_5 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_2022) begin
                              portQ_5 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_2022) begin
                                portQ_5 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_2022) begin
                                  portQ_5 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_2022) begin
                                    portQ_5 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_2022) begin
                                      portQ_5 <= io_bbLoadPorts_1;
                                    end else begin
                                      portQ_5 <= 1'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        if (4'hf == _T_2040) begin
          portQ_6 <= 1'h0;
        end else begin
          if (4'he == _T_2040) begin
            portQ_6 <= 1'h0;
          end else begin
            if (4'hd == _T_2040) begin
              portQ_6 <= 1'h0;
            end else begin
              if (4'hc == _T_2040) begin
                portQ_6 <= 1'h0;
              end else begin
                if (4'hb == _T_2040) begin
                  portQ_6 <= 1'h0;
                end else begin
                  if (4'ha == _T_2040) begin
                    portQ_6 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_2040) begin
                      portQ_6 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_2040) begin
                        portQ_6 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_2040) begin
                          portQ_6 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_2040) begin
                            portQ_6 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_2040) begin
                              portQ_6 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_2040) begin
                                portQ_6 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_2040) begin
                                  portQ_6 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_2040) begin
                                    portQ_6 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_2040) begin
                                      portQ_6 <= io_bbLoadPorts_1;
                                    end else begin
                                      portQ_6 <= 1'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        if (4'hf == _T_2058) begin
          portQ_7 <= 1'h0;
        end else begin
          if (4'he == _T_2058) begin
            portQ_7 <= 1'h0;
          end else begin
            if (4'hd == _T_2058) begin
              portQ_7 <= 1'h0;
            end else begin
              if (4'hc == _T_2058) begin
                portQ_7 <= 1'h0;
              end else begin
                if (4'hb == _T_2058) begin
                  portQ_7 <= 1'h0;
                end else begin
                  if (4'ha == _T_2058) begin
                    portQ_7 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_2058) begin
                      portQ_7 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_2058) begin
                        portQ_7 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_2058) begin
                          portQ_7 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_2058) begin
                            portQ_7 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_2058) begin
                              portQ_7 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_2058) begin
                                portQ_7 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_2058) begin
                                  portQ_7 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_2058) begin
                                    portQ_7 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_2058) begin
                                      portQ_7 <= io_bbLoadPorts_1;
                                    end else begin
                                      portQ_7 <= 1'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        if (4'hf == _T_2076) begin
          portQ_8 <= 1'h0;
        end else begin
          if (4'he == _T_2076) begin
            portQ_8 <= 1'h0;
          end else begin
            if (4'hd == _T_2076) begin
              portQ_8 <= 1'h0;
            end else begin
              if (4'hc == _T_2076) begin
                portQ_8 <= 1'h0;
              end else begin
                if (4'hb == _T_2076) begin
                  portQ_8 <= 1'h0;
                end else begin
                  if (4'ha == _T_2076) begin
                    portQ_8 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_2076) begin
                      portQ_8 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_2076) begin
                        portQ_8 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_2076) begin
                          portQ_8 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_2076) begin
                            portQ_8 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_2076) begin
                              portQ_8 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_2076) begin
                                portQ_8 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_2076) begin
                                  portQ_8 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_2076) begin
                                    portQ_8 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_2076) begin
                                      portQ_8 <= io_bbLoadPorts_1;
                                    end else begin
                                      portQ_8 <= 1'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        if (4'hf == _T_2094) begin
          portQ_9 <= 1'h0;
        end else begin
          if (4'he == _T_2094) begin
            portQ_9 <= 1'h0;
          end else begin
            if (4'hd == _T_2094) begin
              portQ_9 <= 1'h0;
            end else begin
              if (4'hc == _T_2094) begin
                portQ_9 <= 1'h0;
              end else begin
                if (4'hb == _T_2094) begin
                  portQ_9 <= 1'h0;
                end else begin
                  if (4'ha == _T_2094) begin
                    portQ_9 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_2094) begin
                      portQ_9 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_2094) begin
                        portQ_9 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_2094) begin
                          portQ_9 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_2094) begin
                            portQ_9 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_2094) begin
                              portQ_9 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_2094) begin
                                portQ_9 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_2094) begin
                                  portQ_9 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_2094) begin
                                    portQ_9 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_2094) begin
                                      portQ_9 <= io_bbLoadPorts_1;
                                    end else begin
                                      portQ_9 <= 1'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        if (4'hf == _T_2112) begin
          portQ_10 <= 1'h0;
        end else begin
          if (4'he == _T_2112) begin
            portQ_10 <= 1'h0;
          end else begin
            if (4'hd == _T_2112) begin
              portQ_10 <= 1'h0;
            end else begin
              if (4'hc == _T_2112) begin
                portQ_10 <= 1'h0;
              end else begin
                if (4'hb == _T_2112) begin
                  portQ_10 <= 1'h0;
                end else begin
                  if (4'ha == _T_2112) begin
                    portQ_10 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_2112) begin
                      portQ_10 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_2112) begin
                        portQ_10 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_2112) begin
                          portQ_10 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_2112) begin
                            portQ_10 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_2112) begin
                              portQ_10 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_2112) begin
                                portQ_10 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_2112) begin
                                  portQ_10 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_2112) begin
                                    portQ_10 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_2112) begin
                                      portQ_10 <= io_bbLoadPorts_1;
                                    end else begin
                                      portQ_10 <= 1'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        if (4'hf == _T_2130) begin
          portQ_11 <= 1'h0;
        end else begin
          if (4'he == _T_2130) begin
            portQ_11 <= 1'h0;
          end else begin
            if (4'hd == _T_2130) begin
              portQ_11 <= 1'h0;
            end else begin
              if (4'hc == _T_2130) begin
                portQ_11 <= 1'h0;
              end else begin
                if (4'hb == _T_2130) begin
                  portQ_11 <= 1'h0;
                end else begin
                  if (4'ha == _T_2130) begin
                    portQ_11 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_2130) begin
                      portQ_11 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_2130) begin
                        portQ_11 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_2130) begin
                          portQ_11 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_2130) begin
                            portQ_11 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_2130) begin
                              portQ_11 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_2130) begin
                                portQ_11 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_2130) begin
                                  portQ_11 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_2130) begin
                                    portQ_11 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_2130) begin
                                      portQ_11 <= io_bbLoadPorts_1;
                                    end else begin
                                      portQ_11 <= 1'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        if (4'hf == _T_2148) begin
          portQ_12 <= 1'h0;
        end else begin
          if (4'he == _T_2148) begin
            portQ_12 <= 1'h0;
          end else begin
            if (4'hd == _T_2148) begin
              portQ_12 <= 1'h0;
            end else begin
              if (4'hc == _T_2148) begin
                portQ_12 <= 1'h0;
              end else begin
                if (4'hb == _T_2148) begin
                  portQ_12 <= 1'h0;
                end else begin
                  if (4'ha == _T_2148) begin
                    portQ_12 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_2148) begin
                      portQ_12 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_2148) begin
                        portQ_12 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_2148) begin
                          portQ_12 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_2148) begin
                            portQ_12 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_2148) begin
                              portQ_12 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_2148) begin
                                portQ_12 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_2148) begin
                                  portQ_12 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_2148) begin
                                    portQ_12 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_2148) begin
                                      portQ_12 <= io_bbLoadPorts_1;
                                    end else begin
                                      portQ_12 <= 1'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        if (4'hf == _T_2166) begin
          portQ_13 <= 1'h0;
        end else begin
          if (4'he == _T_2166) begin
            portQ_13 <= 1'h0;
          end else begin
            if (4'hd == _T_2166) begin
              portQ_13 <= 1'h0;
            end else begin
              if (4'hc == _T_2166) begin
                portQ_13 <= 1'h0;
              end else begin
                if (4'hb == _T_2166) begin
                  portQ_13 <= 1'h0;
                end else begin
                  if (4'ha == _T_2166) begin
                    portQ_13 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_2166) begin
                      portQ_13 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_2166) begin
                        portQ_13 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_2166) begin
                          portQ_13 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_2166) begin
                            portQ_13 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_2166) begin
                              portQ_13 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_2166) begin
                                portQ_13 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_2166) begin
                                  portQ_13 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_2166) begin
                                    portQ_13 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_2166) begin
                                      portQ_13 <= io_bbLoadPorts_1;
                                    end else begin
                                      portQ_13 <= 1'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        if (4'hf == _T_2184) begin
          portQ_14 <= 1'h0;
        end else begin
          if (4'he == _T_2184) begin
            portQ_14 <= 1'h0;
          end else begin
            if (4'hd == _T_2184) begin
              portQ_14 <= 1'h0;
            end else begin
              if (4'hc == _T_2184) begin
                portQ_14 <= 1'h0;
              end else begin
                if (4'hb == _T_2184) begin
                  portQ_14 <= 1'h0;
                end else begin
                  if (4'ha == _T_2184) begin
                    portQ_14 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_2184) begin
                      portQ_14 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_2184) begin
                        portQ_14 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_2184) begin
                          portQ_14 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_2184) begin
                            portQ_14 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_2184) begin
                              portQ_14 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_2184) begin
                                portQ_14 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_2184) begin
                                  portQ_14 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_2184) begin
                                    portQ_14 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_2184) begin
                                      portQ_14 <= io_bbLoadPorts_1;
                                    end else begin
                                      portQ_14 <= 1'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        if (4'hf == _T_2202) begin
          portQ_15 <= 1'h0;
        end else begin
          if (4'he == _T_2202) begin
            portQ_15 <= 1'h0;
          end else begin
            if (4'hd == _T_2202) begin
              portQ_15 <= 1'h0;
            end else begin
              if (4'hc == _T_2202) begin
                portQ_15 <= 1'h0;
              end else begin
                if (4'hb == _T_2202) begin
                  portQ_15 <= 1'h0;
                end else begin
                  if (4'ha == _T_2202) begin
                    portQ_15 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_2202) begin
                      portQ_15 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_2202) begin
                        portQ_15 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_2202) begin
                          portQ_15 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_2202) begin
                            portQ_15 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_2202) begin
                              portQ_15 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_2202) begin
                                portQ_15 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_2202) begin
                                  portQ_15 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_2202) begin
                                    portQ_15 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_2202) begin
                                      portQ_15 <= io_bbLoadPorts_1;
                                    end else begin
                                      portQ_15 <= 1'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      addrQ_0 <= 32'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_101219) begin
          if (_T_101221) begin
            addrQ_0 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_0 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_1 <= 32'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_101237) begin
          if (_T_101239) begin
            addrQ_1 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_1 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_2 <= 32'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_101255) begin
          if (_T_101257) begin
            addrQ_2 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_2 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_3 <= 32'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_101273) begin
          if (_T_101275) begin
            addrQ_3 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_3 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_4 <= 32'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_101291) begin
          if (_T_101293) begin
            addrQ_4 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_4 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_5 <= 32'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_101309) begin
          if (_T_101311) begin
            addrQ_5 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_5 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_6 <= 32'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_101327) begin
          if (_T_101329) begin
            addrQ_6 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_6 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_7 <= 32'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_101345) begin
          if (_T_101347) begin
            addrQ_7 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_7 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_8 <= 32'h0;
    end else begin
      if (!(initBits_8)) begin
        if (_T_101363) begin
          if (_T_101365) begin
            addrQ_8 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_8 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_9 <= 32'h0;
    end else begin
      if (!(initBits_9)) begin
        if (_T_101381) begin
          if (_T_101383) begin
            addrQ_9 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_9 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_10 <= 32'h0;
    end else begin
      if (!(initBits_10)) begin
        if (_T_101399) begin
          if (_T_101401) begin
            addrQ_10 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_10 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_11 <= 32'h0;
    end else begin
      if (!(initBits_11)) begin
        if (_T_101417) begin
          if (_T_101419) begin
            addrQ_11 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_11 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_12 <= 32'h0;
    end else begin
      if (!(initBits_12)) begin
        if (_T_101435) begin
          if (_T_101437) begin
            addrQ_12 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_12 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_13 <= 32'h0;
    end else begin
      if (!(initBits_13)) begin
        if (_T_101453) begin
          if (_T_101455) begin
            addrQ_13 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_13 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_14 <= 32'h0;
    end else begin
      if (!(initBits_14)) begin
        if (_T_101471) begin
          if (_T_101473) begin
            addrQ_14 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_14 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_15 <= 32'h0;
    end else begin
      if (!(initBits_15)) begin
        if (_T_101489) begin
          if (_T_101491) begin
            addrQ_15 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_15 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_0 <= 32'h0;
    end else begin
      if (bypassRequest_0) begin
        if (_T_88306) begin
          if (4'hf == _T_88289) begin
            dataQ_0 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88289) begin
              dataQ_0 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88289) begin
                dataQ_0 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88289) begin
                  dataQ_0 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88289) begin
                    dataQ_0 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88289) begin
                      dataQ_0 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88289) begin
                        dataQ_0 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88289) begin
                          dataQ_0 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88289) begin
                            dataQ_0 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88289) begin
                              dataQ_0 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88289) begin
                                dataQ_0 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88289) begin
                                  dataQ_0 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88289) begin
                                    dataQ_0 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88289) begin
                                      dataQ_0 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88289) begin
                                        dataQ_0 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_0 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_0 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_0) begin
          dataQ_0 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_1 <= 32'h0;
    end else begin
      if (bypassRequest_1) begin
        if (_T_88442) begin
          if (4'hf == _T_88425) begin
            dataQ_1 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88425) begin
              dataQ_1 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88425) begin
                dataQ_1 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88425) begin
                  dataQ_1 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88425) begin
                    dataQ_1 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88425) begin
                      dataQ_1 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88425) begin
                        dataQ_1 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88425) begin
                          dataQ_1 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88425) begin
                            dataQ_1 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88425) begin
                              dataQ_1 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88425) begin
                                dataQ_1 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88425) begin
                                  dataQ_1 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88425) begin
                                    dataQ_1 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88425) begin
                                      dataQ_1 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88425) begin
                                        dataQ_1 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_1 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_1 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_1) begin
          dataQ_1 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_2 <= 32'h0;
    end else begin
      if (bypassRequest_2) begin
        if (_T_88578) begin
          if (4'hf == _T_88561) begin
            dataQ_2 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88561) begin
              dataQ_2 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88561) begin
                dataQ_2 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88561) begin
                  dataQ_2 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88561) begin
                    dataQ_2 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88561) begin
                      dataQ_2 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88561) begin
                        dataQ_2 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88561) begin
                          dataQ_2 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88561) begin
                            dataQ_2 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88561) begin
                              dataQ_2 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88561) begin
                                dataQ_2 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88561) begin
                                  dataQ_2 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88561) begin
                                    dataQ_2 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88561) begin
                                      dataQ_2 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88561) begin
                                        dataQ_2 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_2 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_2 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_2) begin
          dataQ_2 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_3 <= 32'h0;
    end else begin
      if (bypassRequest_3) begin
        if (_T_88714) begin
          if (4'hf == _T_88697) begin
            dataQ_3 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88697) begin
              dataQ_3 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88697) begin
                dataQ_3 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88697) begin
                  dataQ_3 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88697) begin
                    dataQ_3 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88697) begin
                      dataQ_3 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88697) begin
                        dataQ_3 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88697) begin
                          dataQ_3 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88697) begin
                            dataQ_3 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88697) begin
                              dataQ_3 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88697) begin
                                dataQ_3 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88697) begin
                                  dataQ_3 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88697) begin
                                    dataQ_3 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88697) begin
                                      dataQ_3 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88697) begin
                                        dataQ_3 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_3 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_3 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_3) begin
          dataQ_3 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_4 <= 32'h0;
    end else begin
      if (bypassRequest_4) begin
        if (_T_88850) begin
          if (4'hf == _T_88833) begin
            dataQ_4 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88833) begin
              dataQ_4 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88833) begin
                dataQ_4 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88833) begin
                  dataQ_4 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88833) begin
                    dataQ_4 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88833) begin
                      dataQ_4 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88833) begin
                        dataQ_4 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88833) begin
                          dataQ_4 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88833) begin
                            dataQ_4 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88833) begin
                              dataQ_4 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88833) begin
                                dataQ_4 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88833) begin
                                  dataQ_4 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88833) begin
                                    dataQ_4 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88833) begin
                                      dataQ_4 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88833) begin
                                        dataQ_4 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_4 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_4 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_4) begin
          dataQ_4 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_5 <= 32'h0;
    end else begin
      if (bypassRequest_5) begin
        if (_T_88986) begin
          if (4'hf == _T_88969) begin
            dataQ_5 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88969) begin
              dataQ_5 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88969) begin
                dataQ_5 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88969) begin
                  dataQ_5 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88969) begin
                    dataQ_5 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88969) begin
                      dataQ_5 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88969) begin
                        dataQ_5 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88969) begin
                          dataQ_5 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88969) begin
                            dataQ_5 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88969) begin
                              dataQ_5 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88969) begin
                                dataQ_5 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88969) begin
                                  dataQ_5 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88969) begin
                                    dataQ_5 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88969) begin
                                      dataQ_5 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88969) begin
                                        dataQ_5 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_5 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_5 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_5) begin
          dataQ_5 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_6 <= 32'h0;
    end else begin
      if (bypassRequest_6) begin
        if (_T_89122) begin
          if (4'hf == _T_89105) begin
            dataQ_6 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89105) begin
              dataQ_6 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89105) begin
                dataQ_6 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89105) begin
                  dataQ_6 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89105) begin
                    dataQ_6 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89105) begin
                      dataQ_6 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89105) begin
                        dataQ_6 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89105) begin
                          dataQ_6 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89105) begin
                            dataQ_6 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89105) begin
                              dataQ_6 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89105) begin
                                dataQ_6 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89105) begin
                                  dataQ_6 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89105) begin
                                    dataQ_6 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89105) begin
                                      dataQ_6 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89105) begin
                                        dataQ_6 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_6 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_6 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_6) begin
          dataQ_6 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_7 <= 32'h0;
    end else begin
      if (bypassRequest_7) begin
        if (_T_89258) begin
          if (4'hf == _T_89241) begin
            dataQ_7 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89241) begin
              dataQ_7 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89241) begin
                dataQ_7 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89241) begin
                  dataQ_7 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89241) begin
                    dataQ_7 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89241) begin
                      dataQ_7 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89241) begin
                        dataQ_7 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89241) begin
                          dataQ_7 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89241) begin
                            dataQ_7 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89241) begin
                              dataQ_7 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89241) begin
                                dataQ_7 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89241) begin
                                  dataQ_7 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89241) begin
                                    dataQ_7 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89241) begin
                                      dataQ_7 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89241) begin
                                        dataQ_7 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_7 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_7 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_7) begin
          dataQ_7 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_8 <= 32'h0;
    end else begin
      if (bypassRequest_8) begin
        if (_T_89394) begin
          if (4'hf == _T_89377) begin
            dataQ_8 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89377) begin
              dataQ_8 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89377) begin
                dataQ_8 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89377) begin
                  dataQ_8 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89377) begin
                    dataQ_8 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89377) begin
                      dataQ_8 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89377) begin
                        dataQ_8 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89377) begin
                          dataQ_8 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89377) begin
                            dataQ_8 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89377) begin
                              dataQ_8 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89377) begin
                                dataQ_8 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89377) begin
                                  dataQ_8 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89377) begin
                                    dataQ_8 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89377) begin
                                      dataQ_8 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89377) begin
                                        dataQ_8 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_8 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_8 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_8) begin
          dataQ_8 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_9 <= 32'h0;
    end else begin
      if (bypassRequest_9) begin
        if (_T_89530) begin
          if (4'hf == _T_89513) begin
            dataQ_9 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89513) begin
              dataQ_9 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89513) begin
                dataQ_9 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89513) begin
                  dataQ_9 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89513) begin
                    dataQ_9 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89513) begin
                      dataQ_9 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89513) begin
                        dataQ_9 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89513) begin
                          dataQ_9 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89513) begin
                            dataQ_9 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89513) begin
                              dataQ_9 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89513) begin
                                dataQ_9 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89513) begin
                                  dataQ_9 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89513) begin
                                    dataQ_9 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89513) begin
                                      dataQ_9 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89513) begin
                                        dataQ_9 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_9 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_9 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_9) begin
          dataQ_9 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_10 <= 32'h0;
    end else begin
      if (bypassRequest_10) begin
        if (_T_89666) begin
          if (4'hf == _T_89649) begin
            dataQ_10 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89649) begin
              dataQ_10 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89649) begin
                dataQ_10 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89649) begin
                  dataQ_10 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89649) begin
                    dataQ_10 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89649) begin
                      dataQ_10 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89649) begin
                        dataQ_10 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89649) begin
                          dataQ_10 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89649) begin
                            dataQ_10 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89649) begin
                              dataQ_10 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89649) begin
                                dataQ_10 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89649) begin
                                  dataQ_10 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89649) begin
                                    dataQ_10 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89649) begin
                                      dataQ_10 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89649) begin
                                        dataQ_10 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_10 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_10 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_10) begin
          dataQ_10 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_11 <= 32'h0;
    end else begin
      if (bypassRequest_11) begin
        if (_T_89802) begin
          if (4'hf == _T_89785) begin
            dataQ_11 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89785) begin
              dataQ_11 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89785) begin
                dataQ_11 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89785) begin
                  dataQ_11 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89785) begin
                    dataQ_11 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89785) begin
                      dataQ_11 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89785) begin
                        dataQ_11 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89785) begin
                          dataQ_11 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89785) begin
                            dataQ_11 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89785) begin
                              dataQ_11 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89785) begin
                                dataQ_11 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89785) begin
                                  dataQ_11 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89785) begin
                                    dataQ_11 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89785) begin
                                      dataQ_11 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89785) begin
                                        dataQ_11 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_11 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_11 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_11) begin
          dataQ_11 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_12 <= 32'h0;
    end else begin
      if (bypassRequest_12) begin
        if (_T_89938) begin
          if (4'hf == _T_89921) begin
            dataQ_12 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89921) begin
              dataQ_12 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89921) begin
                dataQ_12 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89921) begin
                  dataQ_12 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89921) begin
                    dataQ_12 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89921) begin
                      dataQ_12 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89921) begin
                        dataQ_12 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89921) begin
                          dataQ_12 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89921) begin
                            dataQ_12 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89921) begin
                              dataQ_12 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89921) begin
                                dataQ_12 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89921) begin
                                  dataQ_12 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89921) begin
                                    dataQ_12 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89921) begin
                                      dataQ_12 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89921) begin
                                        dataQ_12 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_12 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_12 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_12) begin
          dataQ_12 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_13 <= 32'h0;
    end else begin
      if (bypassRequest_13) begin
        if (_T_90074) begin
          if (4'hf == _T_90057) begin
            dataQ_13 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_90057) begin
              dataQ_13 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_90057) begin
                dataQ_13 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_90057) begin
                  dataQ_13 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_90057) begin
                    dataQ_13 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_90057) begin
                      dataQ_13 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_90057) begin
                        dataQ_13 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_90057) begin
                          dataQ_13 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_90057) begin
                            dataQ_13 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_90057) begin
                              dataQ_13 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_90057) begin
                                dataQ_13 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_90057) begin
                                  dataQ_13 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_90057) begin
                                    dataQ_13 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_90057) begin
                                      dataQ_13 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_90057) begin
                                        dataQ_13 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_13 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_13 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_13) begin
          dataQ_13 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_14 <= 32'h0;
    end else begin
      if (bypassRequest_14) begin
        if (_T_90210) begin
          if (4'hf == _T_90193) begin
            dataQ_14 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_90193) begin
              dataQ_14 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_90193) begin
                dataQ_14 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_90193) begin
                  dataQ_14 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_90193) begin
                    dataQ_14 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_90193) begin
                      dataQ_14 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_90193) begin
                        dataQ_14 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_90193) begin
                          dataQ_14 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_90193) begin
                            dataQ_14 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_90193) begin
                              dataQ_14 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_90193) begin
                                dataQ_14 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_90193) begin
                                  dataQ_14 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_90193) begin
                                    dataQ_14 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_90193) begin
                                      dataQ_14 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_90193) begin
                                        dataQ_14 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_14 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_14 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_14) begin
          dataQ_14 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_15 <= 32'h0;
    end else begin
      if (bypassRequest_15) begin
        if (_T_90346) begin
          if (4'hf == _T_90329) begin
            dataQ_15 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_90329) begin
              dataQ_15 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_90329) begin
                dataQ_15 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_90329) begin
                  dataQ_15 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_90329) begin
                    dataQ_15 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_90329) begin
                      dataQ_15 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_90329) begin
                        dataQ_15 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_90329) begin
                          dataQ_15 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_90329) begin
                            dataQ_15 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_90329) begin
                              dataQ_15 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_90329) begin
                                dataQ_15 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_90329) begin
                                  dataQ_15 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_90329) begin
                                    dataQ_15 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_90329) begin
                                      dataQ_15 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_90329) begin
                                        dataQ_15 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_15 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_15 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_15) begin
          dataQ_15 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      addrKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        addrKnown_0 <= 1'h0;
      end else begin
        if (_T_101219) begin
          addrKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        addrKnown_1 <= 1'h0;
      end else begin
        if (_T_101237) begin
          addrKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        addrKnown_2 <= 1'h0;
      end else begin
        if (_T_101255) begin
          addrKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        addrKnown_3 <= 1'h0;
      end else begin
        if (_T_101273) begin
          addrKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        addrKnown_4 <= 1'h0;
      end else begin
        if (_T_101291) begin
          addrKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        addrKnown_5 <= 1'h0;
      end else begin
        if (_T_101309) begin
          addrKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        addrKnown_6 <= 1'h0;
      end else begin
        if (_T_101327) begin
          addrKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        addrKnown_7 <= 1'h0;
      end else begin
        if (_T_101345) begin
          addrKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        addrKnown_8 <= 1'h0;
      end else begin
        if (_T_101363) begin
          addrKnown_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        addrKnown_9 <= 1'h0;
      end else begin
        if (_T_101381) begin
          addrKnown_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        addrKnown_10 <= 1'h0;
      end else begin
        if (_T_101399) begin
          addrKnown_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        addrKnown_11 <= 1'h0;
      end else begin
        if (_T_101417) begin
          addrKnown_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        addrKnown_12 <= 1'h0;
      end else begin
        if (_T_101435) begin
          addrKnown_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        addrKnown_13 <= 1'h0;
      end else begin
        if (_T_101453) begin
          addrKnown_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        addrKnown_14 <= 1'h0;
      end else begin
        if (_T_101471) begin
          addrKnown_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        addrKnown_15 <= 1'h0;
      end else begin
        if (_T_101489) begin
          addrKnown_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        dataKnown_0 <= 1'h0;
      end else begin
        if (_T_93657) begin
          dataKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        dataKnown_1 <= 1'h0;
      end else begin
        if (_T_93660) begin
          dataKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        dataKnown_2 <= 1'h0;
      end else begin
        if (_T_93663) begin
          dataKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        dataKnown_3 <= 1'h0;
      end else begin
        if (_T_93666) begin
          dataKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        dataKnown_4 <= 1'h0;
      end else begin
        if (_T_93669) begin
          dataKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        dataKnown_5 <= 1'h0;
      end else begin
        if (_T_93672) begin
          dataKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        dataKnown_6 <= 1'h0;
      end else begin
        if (_T_93675) begin
          dataKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        dataKnown_7 <= 1'h0;
      end else begin
        if (_T_93678) begin
          dataKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        dataKnown_8 <= 1'h0;
      end else begin
        if (_T_93681) begin
          dataKnown_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        dataKnown_9 <= 1'h0;
      end else begin
        if (_T_93684) begin
          dataKnown_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        dataKnown_10 <= 1'h0;
      end else begin
        if (_T_93687) begin
          dataKnown_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        dataKnown_11 <= 1'h0;
      end else begin
        if (_T_93690) begin
          dataKnown_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        dataKnown_12 <= 1'h0;
      end else begin
        if (_T_93693) begin
          dataKnown_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        dataKnown_13 <= 1'h0;
      end else begin
        if (_T_93696) begin
          dataKnown_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        dataKnown_14 <= 1'h0;
      end else begin
        if (_T_93699) begin
          dataKnown_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        dataKnown_15 <= 1'h0;
      end else begin
        if (_T_93702) begin
          dataKnown_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        loadCompleted_0 <= 1'h0;
      end else begin
        if (loadCompleting_0) begin
          loadCompleted_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        loadCompleted_1 <= 1'h0;
      end else begin
        if (loadCompleting_1) begin
          loadCompleted_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        loadCompleted_2 <= 1'h0;
      end else begin
        if (loadCompleting_2) begin
          loadCompleted_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        loadCompleted_3 <= 1'h0;
      end else begin
        if (loadCompleting_3) begin
          loadCompleted_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        loadCompleted_4 <= 1'h0;
      end else begin
        if (loadCompleting_4) begin
          loadCompleted_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        loadCompleted_5 <= 1'h0;
      end else begin
        if (loadCompleting_5) begin
          loadCompleted_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        loadCompleted_6 <= 1'h0;
      end else begin
        if (loadCompleting_6) begin
          loadCompleted_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        loadCompleted_7 <= 1'h0;
      end else begin
        if (loadCompleting_7) begin
          loadCompleted_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        loadCompleted_8 <= 1'h0;
      end else begin
        if (loadCompleting_8) begin
          loadCompleted_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        loadCompleted_9 <= 1'h0;
      end else begin
        if (loadCompleting_9) begin
          loadCompleted_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        loadCompleted_10 <= 1'h0;
      end else begin
        if (loadCompleting_10) begin
          loadCompleted_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        loadCompleted_11 <= 1'h0;
      end else begin
        if (loadCompleting_11) begin
          loadCompleted_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        loadCompleted_12 <= 1'h0;
      end else begin
        if (loadCompleting_12) begin
          loadCompleted_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        loadCompleted_13 <= 1'h0;
      end else begin
        if (loadCompleting_13) begin
          loadCompleted_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        loadCompleted_14 <= 1'h0;
      end else begin
        if (loadCompleting_14) begin
          loadCompleted_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        loadCompleted_15 <= 1'h0;
      end else begin
        if (loadCompleting_15) begin
          loadCompleted_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      allocatedEntries_0 <= 1'h0;
    end else begin
      allocatedEntries_0 <= _T_1886;
    end
    if (reset) begin
      allocatedEntries_1 <= 1'h0;
    end else begin
      allocatedEntries_1 <= _T_1887;
    end
    if (reset) begin
      allocatedEntries_2 <= 1'h0;
    end else begin
      allocatedEntries_2 <= _T_1888;
    end
    if (reset) begin
      allocatedEntries_3 <= 1'h0;
    end else begin
      allocatedEntries_3 <= _T_1889;
    end
    if (reset) begin
      allocatedEntries_4 <= 1'h0;
    end else begin
      allocatedEntries_4 <= _T_1890;
    end
    if (reset) begin
      allocatedEntries_5 <= 1'h0;
    end else begin
      allocatedEntries_5 <= _T_1891;
    end
    if (reset) begin
      allocatedEntries_6 <= 1'h0;
    end else begin
      allocatedEntries_6 <= _T_1892;
    end
    if (reset) begin
      allocatedEntries_7 <= 1'h0;
    end else begin
      allocatedEntries_7 <= _T_1893;
    end
    if (reset) begin
      allocatedEntries_8 <= 1'h0;
    end else begin
      allocatedEntries_8 <= _T_1894;
    end
    if (reset) begin
      allocatedEntries_9 <= 1'h0;
    end else begin
      allocatedEntries_9 <= _T_1895;
    end
    if (reset) begin
      allocatedEntries_10 <= 1'h0;
    end else begin
      allocatedEntries_10 <= _T_1896;
    end
    if (reset) begin
      allocatedEntries_11 <= 1'h0;
    end else begin
      allocatedEntries_11 <= _T_1897;
    end
    if (reset) begin
      allocatedEntries_12 <= 1'h0;
    end else begin
      allocatedEntries_12 <= _T_1898;
    end
    if (reset) begin
      allocatedEntries_13 <= 1'h0;
    end else begin
      allocatedEntries_13 <= _T_1899;
    end
    if (reset) begin
      allocatedEntries_14 <= 1'h0;
    end else begin
      allocatedEntries_14 <= _T_1900;
    end
    if (reset) begin
      allocatedEntries_15 <= 1'h0;
    end else begin
      allocatedEntries_15 <= _T_1901;
    end
    if (reset) begin
      bypassInitiated_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        bypassInitiated_0 <= 1'h0;
      end else begin
        if (bypassRequest_0) begin
          bypassInitiated_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        bypassInitiated_1 <= 1'h0;
      end else begin
        if (bypassRequest_1) begin
          bypassInitiated_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        bypassInitiated_2 <= 1'h0;
      end else begin
        if (bypassRequest_2) begin
          bypassInitiated_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        bypassInitiated_3 <= 1'h0;
      end else begin
        if (bypassRequest_3) begin
          bypassInitiated_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        bypassInitiated_4 <= 1'h0;
      end else begin
        if (bypassRequest_4) begin
          bypassInitiated_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        bypassInitiated_5 <= 1'h0;
      end else begin
        if (bypassRequest_5) begin
          bypassInitiated_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        bypassInitiated_6 <= 1'h0;
      end else begin
        if (bypassRequest_6) begin
          bypassInitiated_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        bypassInitiated_7 <= 1'h0;
      end else begin
        if (bypassRequest_7) begin
          bypassInitiated_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        bypassInitiated_8 <= 1'h0;
      end else begin
        if (bypassRequest_8) begin
          bypassInitiated_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        bypassInitiated_9 <= 1'h0;
      end else begin
        if (bypassRequest_9) begin
          bypassInitiated_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        bypassInitiated_10 <= 1'h0;
      end else begin
        if (bypassRequest_10) begin
          bypassInitiated_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        bypassInitiated_11 <= 1'h0;
      end else begin
        if (bypassRequest_11) begin
          bypassInitiated_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        bypassInitiated_12 <= 1'h0;
      end else begin
        if (bypassRequest_12) begin
          bypassInitiated_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        bypassInitiated_13 <= 1'h0;
      end else begin
        if (bypassRequest_13) begin
          bypassInitiated_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        bypassInitiated_14 <= 1'h0;
      end else begin
        if (bypassRequest_14) begin
          bypassInitiated_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        bypassInitiated_15 <= 1'h0;
      end else begin
        if (bypassRequest_15) begin
          bypassInitiated_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      checkBits_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        checkBits_0 <= _T_2229;
      end else begin
        if (io_storeEmpty) begin
          checkBits_0 <= 1'h0;
        end else begin
          if (_T_2233) begin
            checkBits_0 <= 1'h0;
          end else begin
            if (_T_2241) begin
              checkBits_0 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        checkBits_1 <= _T_2259;
      end else begin
        if (io_storeEmpty) begin
          checkBits_1 <= 1'h0;
        end else begin
          if (_T_2263) begin
            checkBits_1 <= 1'h0;
          end else begin
            if (_T_2271) begin
              checkBits_1 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        checkBits_2 <= _T_2289;
      end else begin
        if (io_storeEmpty) begin
          checkBits_2 <= 1'h0;
        end else begin
          if (_T_2293) begin
            checkBits_2 <= 1'h0;
          end else begin
            if (_T_2301) begin
              checkBits_2 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        checkBits_3 <= _T_2319;
      end else begin
        if (io_storeEmpty) begin
          checkBits_3 <= 1'h0;
        end else begin
          if (_T_2323) begin
            checkBits_3 <= 1'h0;
          end else begin
            if (_T_2331) begin
              checkBits_3 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        checkBits_4 <= _T_2349;
      end else begin
        if (io_storeEmpty) begin
          checkBits_4 <= 1'h0;
        end else begin
          if (_T_2353) begin
            checkBits_4 <= 1'h0;
          end else begin
            if (_T_2361) begin
              checkBits_4 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        checkBits_5 <= _T_2379;
      end else begin
        if (io_storeEmpty) begin
          checkBits_5 <= 1'h0;
        end else begin
          if (_T_2383) begin
            checkBits_5 <= 1'h0;
          end else begin
            if (_T_2391) begin
              checkBits_5 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        checkBits_6 <= _T_2409;
      end else begin
        if (io_storeEmpty) begin
          checkBits_6 <= 1'h0;
        end else begin
          if (_T_2413) begin
            checkBits_6 <= 1'h0;
          end else begin
            if (_T_2421) begin
              checkBits_6 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        checkBits_7 <= _T_2439;
      end else begin
        if (io_storeEmpty) begin
          checkBits_7 <= 1'h0;
        end else begin
          if (_T_2443) begin
            checkBits_7 <= 1'h0;
          end else begin
            if (_T_2451) begin
              checkBits_7 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        checkBits_8 <= _T_2469;
      end else begin
        if (io_storeEmpty) begin
          checkBits_8 <= 1'h0;
        end else begin
          if (_T_2473) begin
            checkBits_8 <= 1'h0;
          end else begin
            if (_T_2481) begin
              checkBits_8 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        checkBits_9 <= _T_2499;
      end else begin
        if (io_storeEmpty) begin
          checkBits_9 <= 1'h0;
        end else begin
          if (_T_2503) begin
            checkBits_9 <= 1'h0;
          end else begin
            if (_T_2511) begin
              checkBits_9 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        checkBits_10 <= _T_2529;
      end else begin
        if (io_storeEmpty) begin
          checkBits_10 <= 1'h0;
        end else begin
          if (_T_2533) begin
            checkBits_10 <= 1'h0;
          end else begin
            if (_T_2541) begin
              checkBits_10 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        checkBits_11 <= _T_2559;
      end else begin
        if (io_storeEmpty) begin
          checkBits_11 <= 1'h0;
        end else begin
          if (_T_2563) begin
            checkBits_11 <= 1'h0;
          end else begin
            if (_T_2571) begin
              checkBits_11 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        checkBits_12 <= _T_2589;
      end else begin
        if (io_storeEmpty) begin
          checkBits_12 <= 1'h0;
        end else begin
          if (_T_2593) begin
            checkBits_12 <= 1'h0;
          end else begin
            if (_T_2601) begin
              checkBits_12 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        checkBits_13 <= _T_2619;
      end else begin
        if (io_storeEmpty) begin
          checkBits_13 <= 1'h0;
        end else begin
          if (_T_2623) begin
            checkBits_13 <= 1'h0;
          end else begin
            if (_T_2631) begin
              checkBits_13 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        checkBits_14 <= _T_2649;
      end else begin
        if (io_storeEmpty) begin
          checkBits_14 <= 1'h0;
        end else begin
          if (_T_2653) begin
            checkBits_14 <= 1'h0;
          end else begin
            if (_T_2661) begin
              checkBits_14 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        checkBits_15 <= _T_2679;
      end else begin
        if (io_storeEmpty) begin
          checkBits_15 <= 1'h0;
        end else begin
          if (_T_2683) begin
            checkBits_15 <= 1'h0;
          end else begin
            if (_T_2691) begin
              checkBits_15 <= 1'h0;
            end
          end
        end
      end
    end
    previousStoreHead <= io_storeHead;
    conflictPReg_0_0 <= _T_18290[0];
    conflictPReg_0_1 <= _T_18290[1];
    conflictPReg_0_2 <= _T_18290[2];
    conflictPReg_0_3 <= _T_18290[3];
    conflictPReg_0_4 <= _T_18290[4];
    conflictPReg_0_5 <= _T_18290[5];
    conflictPReg_0_6 <= _T_18290[6];
    conflictPReg_0_7 <= _T_18290[7];
    conflictPReg_0_8 <= _T_18290[8];
    conflictPReg_0_9 <= _T_18290[9];
    conflictPReg_0_10 <= _T_18290[10];
    conflictPReg_0_11 <= _T_18290[11];
    conflictPReg_0_12 <= _T_18290[12];
    conflictPReg_0_13 <= _T_18290[13];
    conflictPReg_0_14 <= _T_18290[14];
    conflictPReg_0_15 <= _T_18290[15];
    conflictPReg_1_0 <= _T_19148[0];
    conflictPReg_1_1 <= _T_19148[1];
    conflictPReg_1_2 <= _T_19148[2];
    conflictPReg_1_3 <= _T_19148[3];
    conflictPReg_1_4 <= _T_19148[4];
    conflictPReg_1_5 <= _T_19148[5];
    conflictPReg_1_6 <= _T_19148[6];
    conflictPReg_1_7 <= _T_19148[7];
    conflictPReg_1_8 <= _T_19148[8];
    conflictPReg_1_9 <= _T_19148[9];
    conflictPReg_1_10 <= _T_19148[10];
    conflictPReg_1_11 <= _T_19148[11];
    conflictPReg_1_12 <= _T_19148[12];
    conflictPReg_1_13 <= _T_19148[13];
    conflictPReg_1_14 <= _T_19148[14];
    conflictPReg_1_15 <= _T_19148[15];
    conflictPReg_2_0 <= _T_20006[0];
    conflictPReg_2_1 <= _T_20006[1];
    conflictPReg_2_2 <= _T_20006[2];
    conflictPReg_2_3 <= _T_20006[3];
    conflictPReg_2_4 <= _T_20006[4];
    conflictPReg_2_5 <= _T_20006[5];
    conflictPReg_2_6 <= _T_20006[6];
    conflictPReg_2_7 <= _T_20006[7];
    conflictPReg_2_8 <= _T_20006[8];
    conflictPReg_2_9 <= _T_20006[9];
    conflictPReg_2_10 <= _T_20006[10];
    conflictPReg_2_11 <= _T_20006[11];
    conflictPReg_2_12 <= _T_20006[12];
    conflictPReg_2_13 <= _T_20006[13];
    conflictPReg_2_14 <= _T_20006[14];
    conflictPReg_2_15 <= _T_20006[15];
    conflictPReg_3_0 <= _T_20864[0];
    conflictPReg_3_1 <= _T_20864[1];
    conflictPReg_3_2 <= _T_20864[2];
    conflictPReg_3_3 <= _T_20864[3];
    conflictPReg_3_4 <= _T_20864[4];
    conflictPReg_3_5 <= _T_20864[5];
    conflictPReg_3_6 <= _T_20864[6];
    conflictPReg_3_7 <= _T_20864[7];
    conflictPReg_3_8 <= _T_20864[8];
    conflictPReg_3_9 <= _T_20864[9];
    conflictPReg_3_10 <= _T_20864[10];
    conflictPReg_3_11 <= _T_20864[11];
    conflictPReg_3_12 <= _T_20864[12];
    conflictPReg_3_13 <= _T_20864[13];
    conflictPReg_3_14 <= _T_20864[14];
    conflictPReg_3_15 <= _T_20864[15];
    conflictPReg_4_0 <= _T_21722[0];
    conflictPReg_4_1 <= _T_21722[1];
    conflictPReg_4_2 <= _T_21722[2];
    conflictPReg_4_3 <= _T_21722[3];
    conflictPReg_4_4 <= _T_21722[4];
    conflictPReg_4_5 <= _T_21722[5];
    conflictPReg_4_6 <= _T_21722[6];
    conflictPReg_4_7 <= _T_21722[7];
    conflictPReg_4_8 <= _T_21722[8];
    conflictPReg_4_9 <= _T_21722[9];
    conflictPReg_4_10 <= _T_21722[10];
    conflictPReg_4_11 <= _T_21722[11];
    conflictPReg_4_12 <= _T_21722[12];
    conflictPReg_4_13 <= _T_21722[13];
    conflictPReg_4_14 <= _T_21722[14];
    conflictPReg_4_15 <= _T_21722[15];
    conflictPReg_5_0 <= _T_22580[0];
    conflictPReg_5_1 <= _T_22580[1];
    conflictPReg_5_2 <= _T_22580[2];
    conflictPReg_5_3 <= _T_22580[3];
    conflictPReg_5_4 <= _T_22580[4];
    conflictPReg_5_5 <= _T_22580[5];
    conflictPReg_5_6 <= _T_22580[6];
    conflictPReg_5_7 <= _T_22580[7];
    conflictPReg_5_8 <= _T_22580[8];
    conflictPReg_5_9 <= _T_22580[9];
    conflictPReg_5_10 <= _T_22580[10];
    conflictPReg_5_11 <= _T_22580[11];
    conflictPReg_5_12 <= _T_22580[12];
    conflictPReg_5_13 <= _T_22580[13];
    conflictPReg_5_14 <= _T_22580[14];
    conflictPReg_5_15 <= _T_22580[15];
    conflictPReg_6_0 <= _T_23438[0];
    conflictPReg_6_1 <= _T_23438[1];
    conflictPReg_6_2 <= _T_23438[2];
    conflictPReg_6_3 <= _T_23438[3];
    conflictPReg_6_4 <= _T_23438[4];
    conflictPReg_6_5 <= _T_23438[5];
    conflictPReg_6_6 <= _T_23438[6];
    conflictPReg_6_7 <= _T_23438[7];
    conflictPReg_6_8 <= _T_23438[8];
    conflictPReg_6_9 <= _T_23438[9];
    conflictPReg_6_10 <= _T_23438[10];
    conflictPReg_6_11 <= _T_23438[11];
    conflictPReg_6_12 <= _T_23438[12];
    conflictPReg_6_13 <= _T_23438[13];
    conflictPReg_6_14 <= _T_23438[14];
    conflictPReg_6_15 <= _T_23438[15];
    conflictPReg_7_0 <= _T_24296[0];
    conflictPReg_7_1 <= _T_24296[1];
    conflictPReg_7_2 <= _T_24296[2];
    conflictPReg_7_3 <= _T_24296[3];
    conflictPReg_7_4 <= _T_24296[4];
    conflictPReg_7_5 <= _T_24296[5];
    conflictPReg_7_6 <= _T_24296[6];
    conflictPReg_7_7 <= _T_24296[7];
    conflictPReg_7_8 <= _T_24296[8];
    conflictPReg_7_9 <= _T_24296[9];
    conflictPReg_7_10 <= _T_24296[10];
    conflictPReg_7_11 <= _T_24296[11];
    conflictPReg_7_12 <= _T_24296[12];
    conflictPReg_7_13 <= _T_24296[13];
    conflictPReg_7_14 <= _T_24296[14];
    conflictPReg_7_15 <= _T_24296[15];
    conflictPReg_8_0 <= _T_25154[0];
    conflictPReg_8_1 <= _T_25154[1];
    conflictPReg_8_2 <= _T_25154[2];
    conflictPReg_8_3 <= _T_25154[3];
    conflictPReg_8_4 <= _T_25154[4];
    conflictPReg_8_5 <= _T_25154[5];
    conflictPReg_8_6 <= _T_25154[6];
    conflictPReg_8_7 <= _T_25154[7];
    conflictPReg_8_8 <= _T_25154[8];
    conflictPReg_8_9 <= _T_25154[9];
    conflictPReg_8_10 <= _T_25154[10];
    conflictPReg_8_11 <= _T_25154[11];
    conflictPReg_8_12 <= _T_25154[12];
    conflictPReg_8_13 <= _T_25154[13];
    conflictPReg_8_14 <= _T_25154[14];
    conflictPReg_8_15 <= _T_25154[15];
    conflictPReg_9_0 <= _T_26012[0];
    conflictPReg_9_1 <= _T_26012[1];
    conflictPReg_9_2 <= _T_26012[2];
    conflictPReg_9_3 <= _T_26012[3];
    conflictPReg_9_4 <= _T_26012[4];
    conflictPReg_9_5 <= _T_26012[5];
    conflictPReg_9_6 <= _T_26012[6];
    conflictPReg_9_7 <= _T_26012[7];
    conflictPReg_9_8 <= _T_26012[8];
    conflictPReg_9_9 <= _T_26012[9];
    conflictPReg_9_10 <= _T_26012[10];
    conflictPReg_9_11 <= _T_26012[11];
    conflictPReg_9_12 <= _T_26012[12];
    conflictPReg_9_13 <= _T_26012[13];
    conflictPReg_9_14 <= _T_26012[14];
    conflictPReg_9_15 <= _T_26012[15];
    conflictPReg_10_0 <= _T_26870[0];
    conflictPReg_10_1 <= _T_26870[1];
    conflictPReg_10_2 <= _T_26870[2];
    conflictPReg_10_3 <= _T_26870[3];
    conflictPReg_10_4 <= _T_26870[4];
    conflictPReg_10_5 <= _T_26870[5];
    conflictPReg_10_6 <= _T_26870[6];
    conflictPReg_10_7 <= _T_26870[7];
    conflictPReg_10_8 <= _T_26870[8];
    conflictPReg_10_9 <= _T_26870[9];
    conflictPReg_10_10 <= _T_26870[10];
    conflictPReg_10_11 <= _T_26870[11];
    conflictPReg_10_12 <= _T_26870[12];
    conflictPReg_10_13 <= _T_26870[13];
    conflictPReg_10_14 <= _T_26870[14];
    conflictPReg_10_15 <= _T_26870[15];
    conflictPReg_11_0 <= _T_27728[0];
    conflictPReg_11_1 <= _T_27728[1];
    conflictPReg_11_2 <= _T_27728[2];
    conflictPReg_11_3 <= _T_27728[3];
    conflictPReg_11_4 <= _T_27728[4];
    conflictPReg_11_5 <= _T_27728[5];
    conflictPReg_11_6 <= _T_27728[6];
    conflictPReg_11_7 <= _T_27728[7];
    conflictPReg_11_8 <= _T_27728[8];
    conflictPReg_11_9 <= _T_27728[9];
    conflictPReg_11_10 <= _T_27728[10];
    conflictPReg_11_11 <= _T_27728[11];
    conflictPReg_11_12 <= _T_27728[12];
    conflictPReg_11_13 <= _T_27728[13];
    conflictPReg_11_14 <= _T_27728[14];
    conflictPReg_11_15 <= _T_27728[15];
    conflictPReg_12_0 <= _T_28586[0];
    conflictPReg_12_1 <= _T_28586[1];
    conflictPReg_12_2 <= _T_28586[2];
    conflictPReg_12_3 <= _T_28586[3];
    conflictPReg_12_4 <= _T_28586[4];
    conflictPReg_12_5 <= _T_28586[5];
    conflictPReg_12_6 <= _T_28586[6];
    conflictPReg_12_7 <= _T_28586[7];
    conflictPReg_12_8 <= _T_28586[8];
    conflictPReg_12_9 <= _T_28586[9];
    conflictPReg_12_10 <= _T_28586[10];
    conflictPReg_12_11 <= _T_28586[11];
    conflictPReg_12_12 <= _T_28586[12];
    conflictPReg_12_13 <= _T_28586[13];
    conflictPReg_12_14 <= _T_28586[14];
    conflictPReg_12_15 <= _T_28586[15];
    conflictPReg_13_0 <= _T_29444[0];
    conflictPReg_13_1 <= _T_29444[1];
    conflictPReg_13_2 <= _T_29444[2];
    conflictPReg_13_3 <= _T_29444[3];
    conflictPReg_13_4 <= _T_29444[4];
    conflictPReg_13_5 <= _T_29444[5];
    conflictPReg_13_6 <= _T_29444[6];
    conflictPReg_13_7 <= _T_29444[7];
    conflictPReg_13_8 <= _T_29444[8];
    conflictPReg_13_9 <= _T_29444[9];
    conflictPReg_13_10 <= _T_29444[10];
    conflictPReg_13_11 <= _T_29444[11];
    conflictPReg_13_12 <= _T_29444[12];
    conflictPReg_13_13 <= _T_29444[13];
    conflictPReg_13_14 <= _T_29444[14];
    conflictPReg_13_15 <= _T_29444[15];
    conflictPReg_14_0 <= _T_30302[0];
    conflictPReg_14_1 <= _T_30302[1];
    conflictPReg_14_2 <= _T_30302[2];
    conflictPReg_14_3 <= _T_30302[3];
    conflictPReg_14_4 <= _T_30302[4];
    conflictPReg_14_5 <= _T_30302[5];
    conflictPReg_14_6 <= _T_30302[6];
    conflictPReg_14_7 <= _T_30302[7];
    conflictPReg_14_8 <= _T_30302[8];
    conflictPReg_14_9 <= _T_30302[9];
    conflictPReg_14_10 <= _T_30302[10];
    conflictPReg_14_11 <= _T_30302[11];
    conflictPReg_14_12 <= _T_30302[12];
    conflictPReg_14_13 <= _T_30302[13];
    conflictPReg_14_14 <= _T_30302[14];
    conflictPReg_14_15 <= _T_30302[15];
    conflictPReg_15_0 <= _T_31160[0];
    conflictPReg_15_1 <= _T_31160[1];
    conflictPReg_15_2 <= _T_31160[2];
    conflictPReg_15_3 <= _T_31160[3];
    conflictPReg_15_4 <= _T_31160[4];
    conflictPReg_15_5 <= _T_31160[5];
    conflictPReg_15_6 <= _T_31160[6];
    conflictPReg_15_7 <= _T_31160[7];
    conflictPReg_15_8 <= _T_31160[8];
    conflictPReg_15_9 <= _T_31160[9];
    conflictPReg_15_10 <= _T_31160[10];
    conflictPReg_15_11 <= _T_31160[11];
    conflictPReg_15_12 <= _T_31160[12];
    conflictPReg_15_13 <= _T_31160[13];
    conflictPReg_15_14 <= _T_31160[14];
    conflictPReg_15_15 <= _T_31160[15];
    storeAddrNotKnownFlagsPReg_0_0 <= _T_52614[0];
    storeAddrNotKnownFlagsPReg_0_1 <= _T_52614[1];
    storeAddrNotKnownFlagsPReg_0_2 <= _T_52614[2];
    storeAddrNotKnownFlagsPReg_0_3 <= _T_52614[3];
    storeAddrNotKnownFlagsPReg_0_4 <= _T_52614[4];
    storeAddrNotKnownFlagsPReg_0_5 <= _T_52614[5];
    storeAddrNotKnownFlagsPReg_0_6 <= _T_52614[6];
    storeAddrNotKnownFlagsPReg_0_7 <= _T_52614[7];
    storeAddrNotKnownFlagsPReg_0_8 <= _T_52614[8];
    storeAddrNotKnownFlagsPReg_0_9 <= _T_52614[9];
    storeAddrNotKnownFlagsPReg_0_10 <= _T_52614[10];
    storeAddrNotKnownFlagsPReg_0_11 <= _T_52614[11];
    storeAddrNotKnownFlagsPReg_0_12 <= _T_52614[12];
    storeAddrNotKnownFlagsPReg_0_13 <= _T_52614[13];
    storeAddrNotKnownFlagsPReg_0_14 <= _T_52614[14];
    storeAddrNotKnownFlagsPReg_0_15 <= _T_52614[15];
    storeAddrNotKnownFlagsPReg_1_0 <= _T_53472[0];
    storeAddrNotKnownFlagsPReg_1_1 <= _T_53472[1];
    storeAddrNotKnownFlagsPReg_1_2 <= _T_53472[2];
    storeAddrNotKnownFlagsPReg_1_3 <= _T_53472[3];
    storeAddrNotKnownFlagsPReg_1_4 <= _T_53472[4];
    storeAddrNotKnownFlagsPReg_1_5 <= _T_53472[5];
    storeAddrNotKnownFlagsPReg_1_6 <= _T_53472[6];
    storeAddrNotKnownFlagsPReg_1_7 <= _T_53472[7];
    storeAddrNotKnownFlagsPReg_1_8 <= _T_53472[8];
    storeAddrNotKnownFlagsPReg_1_9 <= _T_53472[9];
    storeAddrNotKnownFlagsPReg_1_10 <= _T_53472[10];
    storeAddrNotKnownFlagsPReg_1_11 <= _T_53472[11];
    storeAddrNotKnownFlagsPReg_1_12 <= _T_53472[12];
    storeAddrNotKnownFlagsPReg_1_13 <= _T_53472[13];
    storeAddrNotKnownFlagsPReg_1_14 <= _T_53472[14];
    storeAddrNotKnownFlagsPReg_1_15 <= _T_53472[15];
    storeAddrNotKnownFlagsPReg_2_0 <= _T_54330[0];
    storeAddrNotKnownFlagsPReg_2_1 <= _T_54330[1];
    storeAddrNotKnownFlagsPReg_2_2 <= _T_54330[2];
    storeAddrNotKnownFlagsPReg_2_3 <= _T_54330[3];
    storeAddrNotKnownFlagsPReg_2_4 <= _T_54330[4];
    storeAddrNotKnownFlagsPReg_2_5 <= _T_54330[5];
    storeAddrNotKnownFlagsPReg_2_6 <= _T_54330[6];
    storeAddrNotKnownFlagsPReg_2_7 <= _T_54330[7];
    storeAddrNotKnownFlagsPReg_2_8 <= _T_54330[8];
    storeAddrNotKnownFlagsPReg_2_9 <= _T_54330[9];
    storeAddrNotKnownFlagsPReg_2_10 <= _T_54330[10];
    storeAddrNotKnownFlagsPReg_2_11 <= _T_54330[11];
    storeAddrNotKnownFlagsPReg_2_12 <= _T_54330[12];
    storeAddrNotKnownFlagsPReg_2_13 <= _T_54330[13];
    storeAddrNotKnownFlagsPReg_2_14 <= _T_54330[14];
    storeAddrNotKnownFlagsPReg_2_15 <= _T_54330[15];
    storeAddrNotKnownFlagsPReg_3_0 <= _T_55188[0];
    storeAddrNotKnownFlagsPReg_3_1 <= _T_55188[1];
    storeAddrNotKnownFlagsPReg_3_2 <= _T_55188[2];
    storeAddrNotKnownFlagsPReg_3_3 <= _T_55188[3];
    storeAddrNotKnownFlagsPReg_3_4 <= _T_55188[4];
    storeAddrNotKnownFlagsPReg_3_5 <= _T_55188[5];
    storeAddrNotKnownFlagsPReg_3_6 <= _T_55188[6];
    storeAddrNotKnownFlagsPReg_3_7 <= _T_55188[7];
    storeAddrNotKnownFlagsPReg_3_8 <= _T_55188[8];
    storeAddrNotKnownFlagsPReg_3_9 <= _T_55188[9];
    storeAddrNotKnownFlagsPReg_3_10 <= _T_55188[10];
    storeAddrNotKnownFlagsPReg_3_11 <= _T_55188[11];
    storeAddrNotKnownFlagsPReg_3_12 <= _T_55188[12];
    storeAddrNotKnownFlagsPReg_3_13 <= _T_55188[13];
    storeAddrNotKnownFlagsPReg_3_14 <= _T_55188[14];
    storeAddrNotKnownFlagsPReg_3_15 <= _T_55188[15];
    storeAddrNotKnownFlagsPReg_4_0 <= _T_56046[0];
    storeAddrNotKnownFlagsPReg_4_1 <= _T_56046[1];
    storeAddrNotKnownFlagsPReg_4_2 <= _T_56046[2];
    storeAddrNotKnownFlagsPReg_4_3 <= _T_56046[3];
    storeAddrNotKnownFlagsPReg_4_4 <= _T_56046[4];
    storeAddrNotKnownFlagsPReg_4_5 <= _T_56046[5];
    storeAddrNotKnownFlagsPReg_4_6 <= _T_56046[6];
    storeAddrNotKnownFlagsPReg_4_7 <= _T_56046[7];
    storeAddrNotKnownFlagsPReg_4_8 <= _T_56046[8];
    storeAddrNotKnownFlagsPReg_4_9 <= _T_56046[9];
    storeAddrNotKnownFlagsPReg_4_10 <= _T_56046[10];
    storeAddrNotKnownFlagsPReg_4_11 <= _T_56046[11];
    storeAddrNotKnownFlagsPReg_4_12 <= _T_56046[12];
    storeAddrNotKnownFlagsPReg_4_13 <= _T_56046[13];
    storeAddrNotKnownFlagsPReg_4_14 <= _T_56046[14];
    storeAddrNotKnownFlagsPReg_4_15 <= _T_56046[15];
    storeAddrNotKnownFlagsPReg_5_0 <= _T_56904[0];
    storeAddrNotKnownFlagsPReg_5_1 <= _T_56904[1];
    storeAddrNotKnownFlagsPReg_5_2 <= _T_56904[2];
    storeAddrNotKnownFlagsPReg_5_3 <= _T_56904[3];
    storeAddrNotKnownFlagsPReg_5_4 <= _T_56904[4];
    storeAddrNotKnownFlagsPReg_5_5 <= _T_56904[5];
    storeAddrNotKnownFlagsPReg_5_6 <= _T_56904[6];
    storeAddrNotKnownFlagsPReg_5_7 <= _T_56904[7];
    storeAddrNotKnownFlagsPReg_5_8 <= _T_56904[8];
    storeAddrNotKnownFlagsPReg_5_9 <= _T_56904[9];
    storeAddrNotKnownFlagsPReg_5_10 <= _T_56904[10];
    storeAddrNotKnownFlagsPReg_5_11 <= _T_56904[11];
    storeAddrNotKnownFlagsPReg_5_12 <= _T_56904[12];
    storeAddrNotKnownFlagsPReg_5_13 <= _T_56904[13];
    storeAddrNotKnownFlagsPReg_5_14 <= _T_56904[14];
    storeAddrNotKnownFlagsPReg_5_15 <= _T_56904[15];
    storeAddrNotKnownFlagsPReg_6_0 <= _T_57762[0];
    storeAddrNotKnownFlagsPReg_6_1 <= _T_57762[1];
    storeAddrNotKnownFlagsPReg_6_2 <= _T_57762[2];
    storeAddrNotKnownFlagsPReg_6_3 <= _T_57762[3];
    storeAddrNotKnownFlagsPReg_6_4 <= _T_57762[4];
    storeAddrNotKnownFlagsPReg_6_5 <= _T_57762[5];
    storeAddrNotKnownFlagsPReg_6_6 <= _T_57762[6];
    storeAddrNotKnownFlagsPReg_6_7 <= _T_57762[7];
    storeAddrNotKnownFlagsPReg_6_8 <= _T_57762[8];
    storeAddrNotKnownFlagsPReg_6_9 <= _T_57762[9];
    storeAddrNotKnownFlagsPReg_6_10 <= _T_57762[10];
    storeAddrNotKnownFlagsPReg_6_11 <= _T_57762[11];
    storeAddrNotKnownFlagsPReg_6_12 <= _T_57762[12];
    storeAddrNotKnownFlagsPReg_6_13 <= _T_57762[13];
    storeAddrNotKnownFlagsPReg_6_14 <= _T_57762[14];
    storeAddrNotKnownFlagsPReg_6_15 <= _T_57762[15];
    storeAddrNotKnownFlagsPReg_7_0 <= _T_58620[0];
    storeAddrNotKnownFlagsPReg_7_1 <= _T_58620[1];
    storeAddrNotKnownFlagsPReg_7_2 <= _T_58620[2];
    storeAddrNotKnownFlagsPReg_7_3 <= _T_58620[3];
    storeAddrNotKnownFlagsPReg_7_4 <= _T_58620[4];
    storeAddrNotKnownFlagsPReg_7_5 <= _T_58620[5];
    storeAddrNotKnownFlagsPReg_7_6 <= _T_58620[6];
    storeAddrNotKnownFlagsPReg_7_7 <= _T_58620[7];
    storeAddrNotKnownFlagsPReg_7_8 <= _T_58620[8];
    storeAddrNotKnownFlagsPReg_7_9 <= _T_58620[9];
    storeAddrNotKnownFlagsPReg_7_10 <= _T_58620[10];
    storeAddrNotKnownFlagsPReg_7_11 <= _T_58620[11];
    storeAddrNotKnownFlagsPReg_7_12 <= _T_58620[12];
    storeAddrNotKnownFlagsPReg_7_13 <= _T_58620[13];
    storeAddrNotKnownFlagsPReg_7_14 <= _T_58620[14];
    storeAddrNotKnownFlagsPReg_7_15 <= _T_58620[15];
    storeAddrNotKnownFlagsPReg_8_0 <= _T_59478[0];
    storeAddrNotKnownFlagsPReg_8_1 <= _T_59478[1];
    storeAddrNotKnownFlagsPReg_8_2 <= _T_59478[2];
    storeAddrNotKnownFlagsPReg_8_3 <= _T_59478[3];
    storeAddrNotKnownFlagsPReg_8_4 <= _T_59478[4];
    storeAddrNotKnownFlagsPReg_8_5 <= _T_59478[5];
    storeAddrNotKnownFlagsPReg_8_6 <= _T_59478[6];
    storeAddrNotKnownFlagsPReg_8_7 <= _T_59478[7];
    storeAddrNotKnownFlagsPReg_8_8 <= _T_59478[8];
    storeAddrNotKnownFlagsPReg_8_9 <= _T_59478[9];
    storeAddrNotKnownFlagsPReg_8_10 <= _T_59478[10];
    storeAddrNotKnownFlagsPReg_8_11 <= _T_59478[11];
    storeAddrNotKnownFlagsPReg_8_12 <= _T_59478[12];
    storeAddrNotKnownFlagsPReg_8_13 <= _T_59478[13];
    storeAddrNotKnownFlagsPReg_8_14 <= _T_59478[14];
    storeAddrNotKnownFlagsPReg_8_15 <= _T_59478[15];
    storeAddrNotKnownFlagsPReg_9_0 <= _T_60336[0];
    storeAddrNotKnownFlagsPReg_9_1 <= _T_60336[1];
    storeAddrNotKnownFlagsPReg_9_2 <= _T_60336[2];
    storeAddrNotKnownFlagsPReg_9_3 <= _T_60336[3];
    storeAddrNotKnownFlagsPReg_9_4 <= _T_60336[4];
    storeAddrNotKnownFlagsPReg_9_5 <= _T_60336[5];
    storeAddrNotKnownFlagsPReg_9_6 <= _T_60336[6];
    storeAddrNotKnownFlagsPReg_9_7 <= _T_60336[7];
    storeAddrNotKnownFlagsPReg_9_8 <= _T_60336[8];
    storeAddrNotKnownFlagsPReg_9_9 <= _T_60336[9];
    storeAddrNotKnownFlagsPReg_9_10 <= _T_60336[10];
    storeAddrNotKnownFlagsPReg_9_11 <= _T_60336[11];
    storeAddrNotKnownFlagsPReg_9_12 <= _T_60336[12];
    storeAddrNotKnownFlagsPReg_9_13 <= _T_60336[13];
    storeAddrNotKnownFlagsPReg_9_14 <= _T_60336[14];
    storeAddrNotKnownFlagsPReg_9_15 <= _T_60336[15];
    storeAddrNotKnownFlagsPReg_10_0 <= _T_61194[0];
    storeAddrNotKnownFlagsPReg_10_1 <= _T_61194[1];
    storeAddrNotKnownFlagsPReg_10_2 <= _T_61194[2];
    storeAddrNotKnownFlagsPReg_10_3 <= _T_61194[3];
    storeAddrNotKnownFlagsPReg_10_4 <= _T_61194[4];
    storeAddrNotKnownFlagsPReg_10_5 <= _T_61194[5];
    storeAddrNotKnownFlagsPReg_10_6 <= _T_61194[6];
    storeAddrNotKnownFlagsPReg_10_7 <= _T_61194[7];
    storeAddrNotKnownFlagsPReg_10_8 <= _T_61194[8];
    storeAddrNotKnownFlagsPReg_10_9 <= _T_61194[9];
    storeAddrNotKnownFlagsPReg_10_10 <= _T_61194[10];
    storeAddrNotKnownFlagsPReg_10_11 <= _T_61194[11];
    storeAddrNotKnownFlagsPReg_10_12 <= _T_61194[12];
    storeAddrNotKnownFlagsPReg_10_13 <= _T_61194[13];
    storeAddrNotKnownFlagsPReg_10_14 <= _T_61194[14];
    storeAddrNotKnownFlagsPReg_10_15 <= _T_61194[15];
    storeAddrNotKnownFlagsPReg_11_0 <= _T_62052[0];
    storeAddrNotKnownFlagsPReg_11_1 <= _T_62052[1];
    storeAddrNotKnownFlagsPReg_11_2 <= _T_62052[2];
    storeAddrNotKnownFlagsPReg_11_3 <= _T_62052[3];
    storeAddrNotKnownFlagsPReg_11_4 <= _T_62052[4];
    storeAddrNotKnownFlagsPReg_11_5 <= _T_62052[5];
    storeAddrNotKnownFlagsPReg_11_6 <= _T_62052[6];
    storeAddrNotKnownFlagsPReg_11_7 <= _T_62052[7];
    storeAddrNotKnownFlagsPReg_11_8 <= _T_62052[8];
    storeAddrNotKnownFlagsPReg_11_9 <= _T_62052[9];
    storeAddrNotKnownFlagsPReg_11_10 <= _T_62052[10];
    storeAddrNotKnownFlagsPReg_11_11 <= _T_62052[11];
    storeAddrNotKnownFlagsPReg_11_12 <= _T_62052[12];
    storeAddrNotKnownFlagsPReg_11_13 <= _T_62052[13];
    storeAddrNotKnownFlagsPReg_11_14 <= _T_62052[14];
    storeAddrNotKnownFlagsPReg_11_15 <= _T_62052[15];
    storeAddrNotKnownFlagsPReg_12_0 <= _T_62910[0];
    storeAddrNotKnownFlagsPReg_12_1 <= _T_62910[1];
    storeAddrNotKnownFlagsPReg_12_2 <= _T_62910[2];
    storeAddrNotKnownFlagsPReg_12_3 <= _T_62910[3];
    storeAddrNotKnownFlagsPReg_12_4 <= _T_62910[4];
    storeAddrNotKnownFlagsPReg_12_5 <= _T_62910[5];
    storeAddrNotKnownFlagsPReg_12_6 <= _T_62910[6];
    storeAddrNotKnownFlagsPReg_12_7 <= _T_62910[7];
    storeAddrNotKnownFlagsPReg_12_8 <= _T_62910[8];
    storeAddrNotKnownFlagsPReg_12_9 <= _T_62910[9];
    storeAddrNotKnownFlagsPReg_12_10 <= _T_62910[10];
    storeAddrNotKnownFlagsPReg_12_11 <= _T_62910[11];
    storeAddrNotKnownFlagsPReg_12_12 <= _T_62910[12];
    storeAddrNotKnownFlagsPReg_12_13 <= _T_62910[13];
    storeAddrNotKnownFlagsPReg_12_14 <= _T_62910[14];
    storeAddrNotKnownFlagsPReg_12_15 <= _T_62910[15];
    storeAddrNotKnownFlagsPReg_13_0 <= _T_63768[0];
    storeAddrNotKnownFlagsPReg_13_1 <= _T_63768[1];
    storeAddrNotKnownFlagsPReg_13_2 <= _T_63768[2];
    storeAddrNotKnownFlagsPReg_13_3 <= _T_63768[3];
    storeAddrNotKnownFlagsPReg_13_4 <= _T_63768[4];
    storeAddrNotKnownFlagsPReg_13_5 <= _T_63768[5];
    storeAddrNotKnownFlagsPReg_13_6 <= _T_63768[6];
    storeAddrNotKnownFlagsPReg_13_7 <= _T_63768[7];
    storeAddrNotKnownFlagsPReg_13_8 <= _T_63768[8];
    storeAddrNotKnownFlagsPReg_13_9 <= _T_63768[9];
    storeAddrNotKnownFlagsPReg_13_10 <= _T_63768[10];
    storeAddrNotKnownFlagsPReg_13_11 <= _T_63768[11];
    storeAddrNotKnownFlagsPReg_13_12 <= _T_63768[12];
    storeAddrNotKnownFlagsPReg_13_13 <= _T_63768[13];
    storeAddrNotKnownFlagsPReg_13_14 <= _T_63768[14];
    storeAddrNotKnownFlagsPReg_13_15 <= _T_63768[15];
    storeAddrNotKnownFlagsPReg_14_0 <= _T_64626[0];
    storeAddrNotKnownFlagsPReg_14_1 <= _T_64626[1];
    storeAddrNotKnownFlagsPReg_14_2 <= _T_64626[2];
    storeAddrNotKnownFlagsPReg_14_3 <= _T_64626[3];
    storeAddrNotKnownFlagsPReg_14_4 <= _T_64626[4];
    storeAddrNotKnownFlagsPReg_14_5 <= _T_64626[5];
    storeAddrNotKnownFlagsPReg_14_6 <= _T_64626[6];
    storeAddrNotKnownFlagsPReg_14_7 <= _T_64626[7];
    storeAddrNotKnownFlagsPReg_14_8 <= _T_64626[8];
    storeAddrNotKnownFlagsPReg_14_9 <= _T_64626[9];
    storeAddrNotKnownFlagsPReg_14_10 <= _T_64626[10];
    storeAddrNotKnownFlagsPReg_14_11 <= _T_64626[11];
    storeAddrNotKnownFlagsPReg_14_12 <= _T_64626[12];
    storeAddrNotKnownFlagsPReg_14_13 <= _T_64626[13];
    storeAddrNotKnownFlagsPReg_14_14 <= _T_64626[14];
    storeAddrNotKnownFlagsPReg_14_15 <= _T_64626[15];
    storeAddrNotKnownFlagsPReg_15_0 <= _T_65484[0];
    storeAddrNotKnownFlagsPReg_15_1 <= _T_65484[1];
    storeAddrNotKnownFlagsPReg_15_2 <= _T_65484[2];
    storeAddrNotKnownFlagsPReg_15_3 <= _T_65484[3];
    storeAddrNotKnownFlagsPReg_15_4 <= _T_65484[4];
    storeAddrNotKnownFlagsPReg_15_5 <= _T_65484[5];
    storeAddrNotKnownFlagsPReg_15_6 <= _T_65484[6];
    storeAddrNotKnownFlagsPReg_15_7 <= _T_65484[7];
    storeAddrNotKnownFlagsPReg_15_8 <= _T_65484[8];
    storeAddrNotKnownFlagsPReg_15_9 <= _T_65484[9];
    storeAddrNotKnownFlagsPReg_15_10 <= _T_65484[10];
    storeAddrNotKnownFlagsPReg_15_11 <= _T_65484[11];
    storeAddrNotKnownFlagsPReg_15_12 <= _T_65484[12];
    storeAddrNotKnownFlagsPReg_15_13 <= _T_65484[13];
    storeAddrNotKnownFlagsPReg_15_14 <= _T_65484[14];
    storeAddrNotKnownFlagsPReg_15_15 <= _T_65484[15];
    shiftedStoreDataKnownPReg_0 <= _T_5980[0];
    shiftedStoreDataKnownPReg_1 <= _T_5980[1];
    shiftedStoreDataKnownPReg_2 <= _T_5980[2];
    shiftedStoreDataKnownPReg_3 <= _T_5980[3];
    shiftedStoreDataKnownPReg_4 <= _T_5980[4];
    shiftedStoreDataKnownPReg_5 <= _T_5980[5];
    shiftedStoreDataKnownPReg_6 <= _T_5980[6];
    shiftedStoreDataKnownPReg_7 <= _T_5980[7];
    shiftedStoreDataKnownPReg_8 <= _T_5980[8];
    shiftedStoreDataKnownPReg_9 <= _T_5980[9];
    shiftedStoreDataKnownPReg_10 <= _T_5980[10];
    shiftedStoreDataKnownPReg_11 <= _T_5980[11];
    shiftedStoreDataKnownPReg_12 <= _T_5980[12];
    shiftedStoreDataKnownPReg_13 <= _T_5980[13];
    shiftedStoreDataKnownPReg_14 <= _T_5980[14];
    shiftedStoreDataKnownPReg_15 <= _T_5980[15];
    shiftedStoreDataQPreg_0 <= _T_5123[31:0];
    shiftedStoreDataQPreg_1 <= _T_5123[63:32];
    shiftedStoreDataQPreg_2 <= _T_5123[95:64];
    shiftedStoreDataQPreg_3 <= _T_5123[127:96];
    shiftedStoreDataQPreg_4 <= _T_5123[159:128];
    shiftedStoreDataQPreg_5 <= _T_5123[191:160];
    shiftedStoreDataQPreg_6 <= _T_5123[223:192];
    shiftedStoreDataQPreg_7 <= _T_5123[255:224];
    shiftedStoreDataQPreg_8 <= _T_5123[287:256];
    shiftedStoreDataQPreg_9 <= _T_5123[319:288];
    shiftedStoreDataQPreg_10 <= _T_5123[351:320];
    shiftedStoreDataQPreg_11 <= _T_5123[383:352];
    shiftedStoreDataQPreg_12 <= _T_5123[415:384];
    shiftedStoreDataQPreg_13 <= _T_5123[447:416];
    shiftedStoreDataQPreg_14 <= _T_5123[479:448];
    shiftedStoreDataQPreg_15 <= _T_5123[511:480];
    addrKnownPReg_0 <= addrKnown_0;
    addrKnownPReg_1 <= addrKnown_1;
    addrKnownPReg_2 <= addrKnown_2;
    addrKnownPReg_3 <= addrKnown_3;
    addrKnownPReg_4 <= addrKnown_4;
    addrKnownPReg_5 <= addrKnown_5;
    addrKnownPReg_6 <= addrKnown_6;
    addrKnownPReg_7 <= addrKnown_7;
    addrKnownPReg_8 <= addrKnown_8;
    addrKnownPReg_9 <= addrKnown_9;
    addrKnownPReg_10 <= addrKnown_10;
    addrKnownPReg_11 <= addrKnown_11;
    addrKnownPReg_12 <= addrKnown_12;
    addrKnownPReg_13 <= addrKnown_13;
    addrKnownPReg_14 <= addrKnown_14;
    addrKnownPReg_15 <= addrKnown_15;
    dataKnownPReg_0 <= dataKnown_0;
    dataKnownPReg_1 <= dataKnown_1;
    dataKnownPReg_2 <= dataKnown_2;
    dataKnownPReg_3 <= dataKnown_3;
    dataKnownPReg_4 <= dataKnown_4;
    dataKnownPReg_5 <= dataKnown_5;
    dataKnownPReg_6 <= dataKnown_6;
    dataKnownPReg_7 <= dataKnown_7;
    dataKnownPReg_8 <= dataKnown_8;
    dataKnownPReg_9 <= dataKnown_9;
    dataKnownPReg_10 <= dataKnown_10;
    dataKnownPReg_11 <= dataKnown_11;
    dataKnownPReg_12 <= dataKnown_12;
    dataKnownPReg_13 <= dataKnown_13;
    dataKnownPReg_14 <= dataKnown_14;
    dataKnownPReg_15 <= dataKnown_15;
    if (reset) begin
      prevPriorityRequest_15 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_15 <= priorityLoadRequest_15;
      end else begin
        prevPriorityRequest_15 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_14 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_14 <= priorityLoadRequest_14;
      end else begin
        prevPriorityRequest_14 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_13 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_13 <= priorityLoadRequest_13;
      end else begin
        prevPriorityRequest_13 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_12 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_12 <= priorityLoadRequest_12;
      end else begin
        prevPriorityRequest_12 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_11 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_11 <= priorityLoadRequest_11;
      end else begin
        prevPriorityRequest_11 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_10 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_10 <= priorityLoadRequest_10;
      end else begin
        prevPriorityRequest_10 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_9 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_9 <= priorityLoadRequest_9;
      end else begin
        prevPriorityRequest_9 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_8 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_8 <= priorityLoadRequest_8;
      end else begin
        prevPriorityRequest_8 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_7 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_7 <= priorityLoadRequest_7;
      end else begin
        prevPriorityRequest_7 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_6 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_6 <= priorityLoadRequest_6;
      end else begin
        prevPriorityRequest_6 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_5 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_5 <= priorityLoadRequest_5;
      end else begin
        prevPriorityRequest_5 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_4 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_4 <= priorityLoadRequest_4;
      end else begin
        prevPriorityRequest_4 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_3 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_3 <= priorityLoadRequest_3;
      end else begin
        prevPriorityRequest_3 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_2 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_2 <= priorityLoadRequest_2;
      end else begin
        prevPriorityRequest_2 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_1 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_1 <= priorityLoadRequest_1;
      end else begin
        prevPriorityRequest_1 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_0 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_0 <= priorityLoadRequest_0;
      end else begin
        prevPriorityRequest_0 <= 1'h0;
      end
    end
  end
endmodule
module GROUP_ALLOCATOR_LSQ_data( // @[:@45084.2]
  output [3:0] io_bbLoadOffsets_0, // @[:@45087.4]
  output [3:0] io_bbLoadOffsets_1, // @[:@45087.4]
  output [3:0] io_bbLoadOffsets_2, // @[:@45087.4]
  output [3:0] io_bbLoadOffsets_3, // @[:@45087.4]
  output [3:0] io_bbLoadOffsets_4, // @[:@45087.4]
  output [3:0] io_bbLoadOffsets_5, // @[:@45087.4]
  output [3:0] io_bbLoadOffsets_6, // @[:@45087.4]
  output [3:0] io_bbLoadOffsets_7, // @[:@45087.4]
  output [3:0] io_bbLoadOffsets_8, // @[:@45087.4]
  output [3:0] io_bbLoadOffsets_9, // @[:@45087.4]
  output [3:0] io_bbLoadOffsets_10, // @[:@45087.4]
  output [3:0] io_bbLoadOffsets_11, // @[:@45087.4]
  output [3:0] io_bbLoadOffsets_12, // @[:@45087.4]
  output [3:0] io_bbLoadOffsets_13, // @[:@45087.4]
  output [3:0] io_bbLoadOffsets_14, // @[:@45087.4]
  output [3:0] io_bbLoadOffsets_15, // @[:@45087.4]
  output       io_bbLoadPorts_1, // @[:@45087.4]
  output [1:0] io_bbNumLoads, // @[:@45087.4]
  input  [3:0] io_loadTail, // @[:@45087.4]
  input  [3:0] io_loadHead, // @[:@45087.4]
  input        io_loadEmpty, // @[:@45087.4]
  output [3:0] io_bbStoreOffsets_0, // @[:@45087.4]
  output [3:0] io_bbStoreOffsets_1, // @[:@45087.4]
  output [3:0] io_bbStoreOffsets_2, // @[:@45087.4]
  output [3:0] io_bbStoreOffsets_3, // @[:@45087.4]
  output [3:0] io_bbStoreOffsets_4, // @[:@45087.4]
  output [3:0] io_bbStoreOffsets_5, // @[:@45087.4]
  output [3:0] io_bbStoreOffsets_6, // @[:@45087.4]
  output [3:0] io_bbStoreOffsets_7, // @[:@45087.4]
  output [3:0] io_bbStoreOffsets_8, // @[:@45087.4]
  output [3:0] io_bbStoreOffsets_9, // @[:@45087.4]
  output [3:0] io_bbStoreOffsets_10, // @[:@45087.4]
  output [3:0] io_bbStoreOffsets_11, // @[:@45087.4]
  output [3:0] io_bbStoreOffsets_12, // @[:@45087.4]
  output [3:0] io_bbStoreOffsets_13, // @[:@45087.4]
  output [3:0] io_bbStoreOffsets_14, // @[:@45087.4]
  output [3:0] io_bbStoreOffsets_15, // @[:@45087.4]
  output       io_bbNumStores, // @[:@45087.4]
  input  [3:0] io_storeTail, // @[:@45087.4]
  input  [3:0] io_storeHead, // @[:@45087.4]
  input        io_storeEmpty, // @[:@45087.4]
  output       io_bbStart, // @[:@45087.4]
  input        io_bbStartSignals_0, // @[:@45087.4]
  input        io_bbStartSignals_1, // @[:@45087.4]
  output       io_readyToPrevious_0, // @[:@45087.4]
  output       io_readyToPrevious_1, // @[:@45087.4]
  output       io_loadPortsEnable_0, // @[:@45087.4]
  output       io_loadPortsEnable_1, // @[:@45087.4]
  output       io_storePortsEnable_0 // @[:@45087.4]
);
  wire  _T_246; // @[GroupAllocator.scala 42:25:@45090.4]
  wire  _T_247; // @[GroupAllocator.scala 42:16:@45091.4]
  wire [4:0] _GEN_68; // @[GroupAllocator.scala 43:36:@45093.6]
  wire [5:0] _T_249; // @[GroupAllocator.scala 43:36:@45093.6]
  wire [5:0] _T_250; // @[GroupAllocator.scala 43:36:@45094.6]
  wire [4:0] _T_251; // @[GroupAllocator.scala 43:36:@45095.6]
  wire [4:0] _GEN_69; // @[GroupAllocator.scala 43:43:@45096.6]
  wire [5:0] _T_252; // @[GroupAllocator.scala 43:43:@45096.6]
  wire [4:0] _T_253; // @[GroupAllocator.scala 43:43:@45097.6]
  wire [4:0] _T_254; // @[GroupAllocator.scala 45:22:@45101.6]
  wire [4:0] _T_255; // @[GroupAllocator.scala 45:22:@45102.6]
  wire [3:0] _T_256; // @[GroupAllocator.scala 45:22:@45103.6]
  wire [4:0] emptyLoadSlots; // @[GroupAllocator.scala 42:34:@45092.4]
  wire  _T_258; // @[GroupAllocator.scala 42:25:@45107.4]
  wire  _T_259; // @[GroupAllocator.scala 42:16:@45108.4]
  wire [4:0] _GEN_70; // @[GroupAllocator.scala 43:36:@45110.6]
  wire [5:0] _T_261; // @[GroupAllocator.scala 43:36:@45110.6]
  wire [5:0] _T_262; // @[GroupAllocator.scala 43:36:@45111.6]
  wire [4:0] _T_263; // @[GroupAllocator.scala 43:36:@45112.6]
  wire [4:0] _GEN_71; // @[GroupAllocator.scala 43:43:@45113.6]
  wire [5:0] _T_264; // @[GroupAllocator.scala 43:43:@45113.6]
  wire [4:0] _T_265; // @[GroupAllocator.scala 43:43:@45114.6]
  wire [4:0] _T_266; // @[GroupAllocator.scala 45:22:@45118.6]
  wire [4:0] _T_267; // @[GroupAllocator.scala 45:22:@45119.6]
  wire [3:0] _T_268; // @[GroupAllocator.scala 45:22:@45120.6]
  wire [4:0] emptyStoreSlots; // @[GroupAllocator.scala 42:34:@45109.4]
  wire  possibleAllocations_0; // @[GroupAllocator.scala 56:106:@45134.4]
  wire  possibleAllocations_1; // @[GroupAllocator.scala 56:106:@45135.4]
  wire  allocatedBBIdx; // @[Mux.scala 31:69:@45139.4]
  wire  _T_308; // @[GroupAllocator.scala 78:44:@45149.4]
  wire [1:0] _T_470; // @[Mux.scala 46:16:@45288.6]
  wire [1:0] _T_472; // @[Mux.scala 46:16:@45290.6]
  wire  _T_636_1; // @[Mux.scala 46:16:@45351.6]
  wire [5:0] _T_903; // @[GroupAllocator.scala 110:34:@45456.6]
  wire [4:0] _T_904; // @[GroupAllocator.scala 110:34:@45457.6]
  wire [5:0] _T_906; // @[GroupAllocator.scala 110:55:@45458.6]
  wire [5:0] _T_907; // @[GroupAllocator.scala 110:55:@45459.6]
  wire [4:0] _T_908; // @[GroupAllocator.scala 110:55:@45460.6]
  wire [5:0] _T_910; // @[util.scala 10:8:@45461.6]
  wire [5:0] _GEN_0; // @[util.scala 10:14:@45462.6]
  wire [4:0] _T_911; // @[util.scala 10:14:@45462.6]
  wire [3:0] _T_1161; // @[GroupAllocator.scala 110:90:@45624.6 GroupAllocator.scala 110:90:@45625.6]
  wire [3:0] _T_1395_0; // @[Mux.scala 46:16:@45779.6]
  wire [3:0] _T_1432_0; // @[Mux.scala 46:16:@45781.6]
  wire [5:0] _T_1509; // @[GroupAllocator.scala 115:33:@45815.6]
  wire [4:0] _T_1510; // @[GroupAllocator.scala 115:33:@45816.6]
  wire [5:0] _T_1512; // @[GroupAllocator.scala 115:54:@45817.6]
  wire [5:0] _T_1513; // @[GroupAllocator.scala 115:54:@45818.6]
  wire [4:0] _T_1514; // @[GroupAllocator.scala 115:54:@45819.6]
  wire [5:0] _T_1516; // @[util.scala 10:8:@45820.6]
  wire [5:0] _GEN_1; // @[util.scala 10:14:@45821.6]
  wire [4:0] _T_1517; // @[util.scala 10:14:@45821.6]
  wire [3:0] _T_1767; // @[GroupAllocator.scala 115:89:@45983.6 GroupAllocator.scala 115:89:@45984.6]
  wire [3:0] _T_2001_0; // @[Mux.scala 46:16:@46138.6]
  wire [3:0] _T_2038_0; // @[Mux.scala 46:16:@46140.6]
  assign _T_246 = io_loadHead < io_loadTail; // @[GroupAllocator.scala 42:25:@45090.4]
  assign _T_247 = io_loadEmpty | _T_246; // @[GroupAllocator.scala 42:16:@45091.4]
  assign _GEN_68 = {{1'd0}, io_loadTail}; // @[GroupAllocator.scala 43:36:@45093.6]
  assign _T_249 = 5'h10 - _GEN_68; // @[GroupAllocator.scala 43:36:@45093.6]
  assign _T_250 = $unsigned(_T_249); // @[GroupAllocator.scala 43:36:@45094.6]
  assign _T_251 = _T_250[4:0]; // @[GroupAllocator.scala 43:36:@45095.6]
  assign _GEN_69 = {{1'd0}, io_loadHead}; // @[GroupAllocator.scala 43:43:@45096.6]
  assign _T_252 = _T_251 + _GEN_69; // @[GroupAllocator.scala 43:43:@45096.6]
  assign _T_253 = _T_251 + _GEN_69; // @[GroupAllocator.scala 43:43:@45097.6]
  assign _T_254 = io_loadHead - io_loadTail; // @[GroupAllocator.scala 45:22:@45101.6]
  assign _T_255 = $unsigned(_T_254); // @[GroupAllocator.scala 45:22:@45102.6]
  assign _T_256 = _T_255[3:0]; // @[GroupAllocator.scala 45:22:@45103.6]
  assign emptyLoadSlots = _T_247 ? _T_253 : {{1'd0}, _T_256}; // @[GroupAllocator.scala 42:34:@45092.4]
  assign _T_258 = io_storeHead < io_storeTail; // @[GroupAllocator.scala 42:25:@45107.4]
  assign _T_259 = io_storeEmpty | _T_258; // @[GroupAllocator.scala 42:16:@45108.4]
  assign _GEN_70 = {{1'd0}, io_storeTail}; // @[GroupAllocator.scala 43:36:@45110.6]
  assign _T_261 = 5'h10 - _GEN_70; // @[GroupAllocator.scala 43:36:@45110.6]
  assign _T_262 = $unsigned(_T_261); // @[GroupAllocator.scala 43:36:@45111.6]
  assign _T_263 = _T_262[4:0]; // @[GroupAllocator.scala 43:36:@45112.6]
  assign _GEN_71 = {{1'd0}, io_storeHead}; // @[GroupAllocator.scala 43:43:@45113.6]
  assign _T_264 = _T_263 + _GEN_71; // @[GroupAllocator.scala 43:43:@45113.6]
  assign _T_265 = _T_263 + _GEN_71; // @[GroupAllocator.scala 43:43:@45114.6]
  assign _T_266 = io_storeHead - io_storeTail; // @[GroupAllocator.scala 45:22:@45118.6]
  assign _T_267 = $unsigned(_T_266); // @[GroupAllocator.scala 45:22:@45119.6]
  assign _T_268 = _T_267[3:0]; // @[GroupAllocator.scala 45:22:@45120.6]
  assign emptyStoreSlots = _T_259 ? _T_265 : {{1'd0}, _T_268}; // @[GroupAllocator.scala 42:34:@45109.4]
  assign possibleAllocations_0 = io_readyToPrevious_0 & io_bbStartSignals_0; // @[GroupAllocator.scala 56:106:@45134.4]
  assign possibleAllocations_1 = io_readyToPrevious_1 & io_bbStartSignals_1; // @[GroupAllocator.scala 56:106:@45135.4]
  assign allocatedBBIdx = possibleAllocations_0 ? 1'h0 : 1'h1; // @[Mux.scala 31:69:@45139.4]
  assign _T_308 = 1'h0 == allocatedBBIdx; // @[GroupAllocator.scala 78:44:@45149.4]
  assign _T_470 = allocatedBBIdx ? 2'h2 : 2'h0; // @[Mux.scala 46:16:@45288.6]
  assign _T_472 = _T_308 ? 2'h0 : _T_470; // @[Mux.scala 46:16:@45290.6]
  assign _T_636_1 = _T_308 ? 1'h0 : allocatedBBIdx; // @[Mux.scala 46:16:@45351.6]
  assign _T_903 = _GEN_70 + 5'h10; // @[GroupAllocator.scala 110:34:@45456.6]
  assign _T_904 = _GEN_70 + 5'h10; // @[GroupAllocator.scala 110:34:@45457.6]
  assign _T_906 = _T_904 - 5'h1; // @[GroupAllocator.scala 110:55:@45458.6]
  assign _T_907 = $unsigned(_T_906); // @[GroupAllocator.scala 110:55:@45459.6]
  assign _T_908 = _T_907[4:0]; // @[GroupAllocator.scala 110:55:@45460.6]
  assign _T_910 = {{1'd0}, _T_908}; // @[util.scala 10:8:@45461.6]
  assign _GEN_0 = _T_910 % 6'h10; // @[util.scala 10:14:@45462.6]
  assign _T_911 = _GEN_0[4:0]; // @[util.scala 10:14:@45462.6]
  assign _T_1161 = _T_911[3:0]; // @[GroupAllocator.scala 110:90:@45624.6 GroupAllocator.scala 110:90:@45625.6]
  assign _T_1395_0 = allocatedBBIdx ? _T_1161 : 4'h0; // @[Mux.scala 46:16:@45779.6]
  assign _T_1432_0 = _T_308 ? _T_1161 : _T_1395_0; // @[Mux.scala 46:16:@45781.6]
  assign _T_1509 = _GEN_68 + 5'h10; // @[GroupAllocator.scala 115:33:@45815.6]
  assign _T_1510 = _GEN_68 + 5'h10; // @[GroupAllocator.scala 115:33:@45816.6]
  assign _T_1512 = _T_1510 - 5'h1; // @[GroupAllocator.scala 115:54:@45817.6]
  assign _T_1513 = $unsigned(_T_1512); // @[GroupAllocator.scala 115:54:@45818.6]
  assign _T_1514 = _T_1513[4:0]; // @[GroupAllocator.scala 115:54:@45819.6]
  assign _T_1516 = {{1'd0}, _T_1514}; // @[util.scala 10:8:@45820.6]
  assign _GEN_1 = _T_1516 % 6'h10; // @[util.scala 10:14:@45821.6]
  assign _T_1517 = _GEN_1[4:0]; // @[util.scala 10:14:@45821.6]
  assign _T_1767 = _T_1517[3:0]; // @[GroupAllocator.scala 115:89:@45983.6 GroupAllocator.scala 115:89:@45984.6]
  assign _T_2001_0 = allocatedBBIdx ? _T_1767 : 4'h0; // @[Mux.scala 46:16:@46138.6]
  assign _T_2038_0 = _T_308 ? _T_1767 : _T_2001_0; // @[Mux.scala 46:16:@46140.6]
  assign io_bbLoadOffsets_0 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45237.4 GroupAllocator.scala 106:22:@45782.6]
  assign io_bbLoadOffsets_1 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45238.4 GroupAllocator.scala 106:22:@45783.6]
  assign io_bbLoadOffsets_2 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45239.4 GroupAllocator.scala 106:22:@45784.6]
  assign io_bbLoadOffsets_3 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45240.4 GroupAllocator.scala 106:22:@45785.6]
  assign io_bbLoadOffsets_4 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45241.4 GroupAllocator.scala 106:22:@45786.6]
  assign io_bbLoadOffsets_5 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45242.4 GroupAllocator.scala 106:22:@45787.6]
  assign io_bbLoadOffsets_6 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45243.4 GroupAllocator.scala 106:22:@45788.6]
  assign io_bbLoadOffsets_7 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45244.4 GroupAllocator.scala 106:22:@45789.6]
  assign io_bbLoadOffsets_8 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45245.4 GroupAllocator.scala 106:22:@45790.6]
  assign io_bbLoadOffsets_9 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45246.4 GroupAllocator.scala 106:22:@45791.6]
  assign io_bbLoadOffsets_10 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45247.4 GroupAllocator.scala 106:22:@45792.6]
  assign io_bbLoadOffsets_11 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45248.4 GroupAllocator.scala 106:22:@45793.6]
  assign io_bbLoadOffsets_12 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45249.4 GroupAllocator.scala 106:22:@45794.6]
  assign io_bbLoadOffsets_13 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45250.4 GroupAllocator.scala 106:22:@45795.6]
  assign io_bbLoadOffsets_14 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45251.4 GroupAllocator.scala 106:22:@45796.6]
  assign io_bbLoadOffsets_15 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45252.4 GroupAllocator.scala 106:22:@45797.6]
  assign io_bbLoadPorts_1 = io_bbStart ? _T_636_1 : 1'h0; // @[GroupAllocator.scala 87:18:@45172.4 GroupAllocator.scala 95:20:@45353.6]
  assign io_bbNumLoads = io_bbStart ? _T_472 : 2'h0; // @[GroupAllocator.scala 85:17:@45152.4 GroupAllocator.scala 93:19:@45291.6]
  assign io_bbStoreOffsets_0 = io_bbStart ? _T_2038_0 : 4'h0; // @[GroupAllocator.scala 90:21:@45270.4 GroupAllocator.scala 111:23:@46141.6]
  assign io_bbStoreOffsets_1 = io_bbStart ? _T_2038_0 : 4'h0; // @[GroupAllocator.scala 90:21:@45271.4 GroupAllocator.scala 111:23:@46142.6]
  assign io_bbStoreOffsets_2 = io_bbStart ? _T_2038_0 : 4'h0; // @[GroupAllocator.scala 90:21:@45272.4 GroupAllocator.scala 111:23:@46143.6]
  assign io_bbStoreOffsets_3 = io_bbStart ? _T_2038_0 : 4'h0; // @[GroupAllocator.scala 90:21:@45273.4 GroupAllocator.scala 111:23:@46144.6]
  assign io_bbStoreOffsets_4 = io_bbStart ? _T_2038_0 : 4'h0; // @[GroupAllocator.scala 90:21:@45274.4 GroupAllocator.scala 111:23:@46145.6]
  assign io_bbStoreOffsets_5 = io_bbStart ? _T_2038_0 : 4'h0; // @[GroupAllocator.scala 90:21:@45275.4 GroupAllocator.scala 111:23:@46146.6]
  assign io_bbStoreOffsets_6 = io_bbStart ? _T_2038_0 : 4'h0; // @[GroupAllocator.scala 90:21:@45276.4 GroupAllocator.scala 111:23:@46147.6]
  assign io_bbStoreOffsets_7 = io_bbStart ? _T_2038_0 : 4'h0; // @[GroupAllocator.scala 90:21:@45277.4 GroupAllocator.scala 111:23:@46148.6]
  assign io_bbStoreOffsets_8 = io_bbStart ? _T_2038_0 : 4'h0; // @[GroupAllocator.scala 90:21:@45278.4 GroupAllocator.scala 111:23:@46149.6]
  assign io_bbStoreOffsets_9 = io_bbStart ? _T_2038_0 : 4'h0; // @[GroupAllocator.scala 90:21:@45279.4 GroupAllocator.scala 111:23:@46150.6]
  assign io_bbStoreOffsets_10 = io_bbStart ? _T_2038_0 : 4'h0; // @[GroupAllocator.scala 90:21:@45280.4 GroupAllocator.scala 111:23:@46151.6]
  assign io_bbStoreOffsets_11 = io_bbStart ? _T_2038_0 : 4'h0; // @[GroupAllocator.scala 90:21:@45281.4 GroupAllocator.scala 111:23:@46152.6]
  assign io_bbStoreOffsets_12 = io_bbStart ? _T_2038_0 : 4'h0; // @[GroupAllocator.scala 90:21:@45282.4 GroupAllocator.scala 111:23:@46153.6]
  assign io_bbStoreOffsets_13 = io_bbStart ? _T_2038_0 : 4'h0; // @[GroupAllocator.scala 90:21:@45283.4 GroupAllocator.scala 111:23:@46154.6]
  assign io_bbStoreOffsets_14 = io_bbStart ? _T_2038_0 : 4'h0; // @[GroupAllocator.scala 90:21:@45284.4 GroupAllocator.scala 111:23:@46155.6]
  assign io_bbStoreOffsets_15 = io_bbStart ? _T_2038_0 : 4'h0; // @[GroupAllocator.scala 90:21:@45285.4 GroupAllocator.scala 111:23:@46156.6]
  assign io_bbNumStores = io_bbStart ? _T_308 : 1'h0; // @[GroupAllocator.scala 86:18:@45153.4 GroupAllocator.scala 94:20:@45296.6]
  assign io_bbStart = possibleAllocations_0 | possibleAllocations_1; // @[GroupAllocator.scala 59:14:@45142.4]
  assign io_readyToPrevious_0 = 5'h1 <= emptyStoreSlots; // @[GroupAllocator.scala 53:22:@45132.4]
  assign io_readyToPrevious_1 = 5'h2 <= emptyLoadSlots; // @[GroupAllocator.scala 53:22:@45133.4]
  assign io_loadPortsEnable_0 = allocatedBBIdx & io_bbStart; // @[GroupAllocator.scala 69:29:@45145.4]
  assign io_loadPortsEnable_1 = allocatedBBIdx & io_bbStart; // @[GroupAllocator.scala 69:29:@45148.4]
  assign io_storePortsEnable_0 = _T_308 & io_bbStart; // @[GroupAllocator.scala 78:30:@45151.4]
endmodule
module LOAD_PORT_LSQ_data( // @[:@46159.2]
  input         clock, // @[:@46160.4]
  input         reset, // @[:@46161.4]
  output        io_addrFromPrev_ready, // @[:@46162.4]
  input         io_addrFromPrev_valid, // @[:@46162.4]
  input  [31:0] io_addrFromPrev_bits, // @[:@46162.4]
  input         io_portEnable, // @[:@46162.4]
  input         io_dataToNext_ready, // @[:@46162.4]
  output        io_dataToNext_valid, // @[:@46162.4]
  output [31:0] io_dataToNext_bits, // @[:@46162.4]
  output        io_loadAddrEnable, // @[:@46162.4]
  output [31:0] io_addrToLoadQueue, // @[:@46162.4]
  output        io_dataFromLoadQueue_ready, // @[:@46162.4]
  input         io_dataFromLoadQueue_valid, // @[:@46162.4]
  input  [31:0] io_dataFromLoadQueue_bits // @[:@46162.4]
);
  reg [4:0] cnt; // @[LoadPort.scala 23:20:@46164.4]
  reg [31:0] _RAND_0;
  wire  _T_44; // @[LoadPort.scala 26:25:@46165.4]
  wire  _T_45; // @[LoadPort.scala 26:22:@46166.4]
  wire  _T_47; // @[LoadPort.scala 26:51:@46167.4]
  wire  _T_48; // @[LoadPort.scala 26:44:@46168.4]
  wire [5:0] _T_50; // @[LoadPort.scala 27:16:@46170.6]
  wire [4:0] _T_51; // @[LoadPort.scala 27:16:@46171.6]
  wire  _T_53; // @[LoadPort.scala 28:35:@46175.6]
  wire  _T_54; // @[LoadPort.scala 28:32:@46176.6]
  wire  _T_56; // @[LoadPort.scala 28:57:@46177.6]
  wire  _T_57; // @[LoadPort.scala 28:50:@46178.6]
  wire [5:0] _T_59; // @[LoadPort.scala 29:16:@46180.8]
  wire [5:0] _T_60; // @[LoadPort.scala 29:16:@46181.8]
  wire [4:0] _T_61; // @[LoadPort.scala 29:16:@46182.8]
  wire [4:0] _GEN_0; // @[LoadPort.scala 28:66:@46179.6]
  wire [4:0] _GEN_1; // @[LoadPort.scala 26:75:@46169.4]
  wire  _T_63; // @[LoadPort.scala 33:28:@46186.4]
  assign _T_44 = io_loadAddrEnable == 1'h0; // @[LoadPort.scala 26:25:@46165.4]
  assign _T_45 = io_portEnable & _T_44; // @[LoadPort.scala 26:22:@46166.4]
  assign _T_47 = cnt != 5'h10; // @[LoadPort.scala 26:51:@46167.4]
  assign _T_48 = _T_45 & _T_47; // @[LoadPort.scala 26:44:@46168.4]
  assign _T_50 = cnt + 5'h1; // @[LoadPort.scala 27:16:@46170.6]
  assign _T_51 = cnt + 5'h1; // @[LoadPort.scala 27:16:@46171.6]
  assign _T_53 = io_portEnable == 1'h0; // @[LoadPort.scala 28:35:@46175.6]
  assign _T_54 = io_loadAddrEnable & _T_53; // @[LoadPort.scala 28:32:@46176.6]
  assign _T_56 = cnt != 5'h0; // @[LoadPort.scala 28:57:@46177.6]
  assign _T_57 = _T_54 & _T_56; // @[LoadPort.scala 28:50:@46178.6]
  assign _T_59 = cnt - 5'h1; // @[LoadPort.scala 29:16:@46180.8]
  assign _T_60 = $unsigned(_T_59); // @[LoadPort.scala 29:16:@46181.8]
  assign _T_61 = _T_60[4:0]; // @[LoadPort.scala 29:16:@46182.8]
  assign _GEN_0 = _T_57 ? _T_61 : cnt; // @[LoadPort.scala 28:66:@46179.6]
  assign _GEN_1 = _T_48 ? _T_51 : _GEN_0; // @[LoadPort.scala 26:75:@46169.4]
  assign _T_63 = cnt > 5'h0; // @[LoadPort.scala 33:28:@46186.4]
  assign io_addrFromPrev_ready = cnt > 5'h0; // @[LoadPort.scala 34:25:@46190.4]
  assign io_dataToNext_valid = io_dataFromLoadQueue_valid; // @[LoadPort.scala 35:17:@46192.4]
  assign io_dataToNext_bits = io_dataFromLoadQueue_bits; // @[LoadPort.scala 35:17:@46191.4]
  assign io_loadAddrEnable = _T_63 & io_addrFromPrev_valid; // @[LoadPort.scala 33:21:@46188.4]
  assign io_addrToLoadQueue = io_addrFromPrev_bits; // @[LoadPort.scala 32:22:@46185.4]
  assign io_dataFromLoadQueue_ready = io_dataToNext_ready; // @[LoadPort.scala 35:17:@46193.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 5'h0;
    end else begin
      if (_T_48) begin
        cnt <= _T_51;
      end else begin
        if (_T_57) begin
          cnt <= _T_61;
        end
      end
    end
  end
endmodule
module STORE_DATA_PORT_LSQ_data( // @[:@46231.2]
  input         clock, // @[:@46232.4]
  input         reset, // @[:@46233.4]
  output        io_dataFromPrev_ready, // @[:@46234.4]
  input         io_dataFromPrev_valid, // @[:@46234.4]
  input  [31:0] io_dataFromPrev_bits, // @[:@46234.4]
  input         io_portEnable, // @[:@46234.4]
  output        io_storeDataEnable, // @[:@46234.4]
  output [31:0] io_dataToStoreQueue // @[:@46234.4]
);
  reg [4:0] cnt; // @[StoreDataPort.scala 21:20:@46236.4]
  reg [31:0] _RAND_0;
  wire  _T_26; // @[StoreDataPort.scala 24:25:@46237.4]
  wire  _T_27; // @[StoreDataPort.scala 24:22:@46238.4]
  wire  _T_29; // @[StoreDataPort.scala 24:52:@46239.4]
  wire  _T_30; // @[StoreDataPort.scala 24:45:@46240.4]
  wire [5:0] _T_32; // @[StoreDataPort.scala 25:16:@46242.6]
  wire [4:0] _T_33; // @[StoreDataPort.scala 25:16:@46243.6]
  wire  _T_35; // @[StoreDataPort.scala 26:36:@46247.6]
  wire  _T_36; // @[StoreDataPort.scala 26:33:@46248.6]
  wire  _T_38; // @[StoreDataPort.scala 26:58:@46249.6]
  wire  _T_39; // @[StoreDataPort.scala 26:51:@46250.6]
  wire [5:0] _T_41; // @[StoreDataPort.scala 27:16:@46252.8]
  wire [5:0] _T_42; // @[StoreDataPort.scala 27:16:@46253.8]
  wire [4:0] _T_43; // @[StoreDataPort.scala 27:16:@46254.8]
  wire [4:0] _GEN_0; // @[StoreDataPort.scala 26:67:@46251.6]
  wire [4:0] _GEN_1; // @[StoreDataPort.scala 24:76:@46241.4]
  wire  _T_45; // @[StoreDataPort.scala 31:29:@46258.4]
  assign _T_26 = io_storeDataEnable == 1'h0; // @[StoreDataPort.scala 24:25:@46237.4]
  assign _T_27 = io_portEnable & _T_26; // @[StoreDataPort.scala 24:22:@46238.4]
  assign _T_29 = cnt != 5'h10; // @[StoreDataPort.scala 24:52:@46239.4]
  assign _T_30 = _T_27 & _T_29; // @[StoreDataPort.scala 24:45:@46240.4]
  assign _T_32 = cnt + 5'h1; // @[StoreDataPort.scala 25:16:@46242.6]
  assign _T_33 = cnt + 5'h1; // @[StoreDataPort.scala 25:16:@46243.6]
  assign _T_35 = io_portEnable == 1'h0; // @[StoreDataPort.scala 26:36:@46247.6]
  assign _T_36 = io_storeDataEnable & _T_35; // @[StoreDataPort.scala 26:33:@46248.6]
  assign _T_38 = cnt != 5'h0; // @[StoreDataPort.scala 26:58:@46249.6]
  assign _T_39 = _T_36 & _T_38; // @[StoreDataPort.scala 26:51:@46250.6]
  assign _T_41 = cnt - 5'h1; // @[StoreDataPort.scala 27:16:@46252.8]
  assign _T_42 = $unsigned(_T_41); // @[StoreDataPort.scala 27:16:@46253.8]
  assign _T_43 = _T_42[4:0]; // @[StoreDataPort.scala 27:16:@46254.8]
  assign _GEN_0 = _T_39 ? _T_43 : cnt; // @[StoreDataPort.scala 26:67:@46251.6]
  assign _GEN_1 = _T_30 ? _T_33 : _GEN_0; // @[StoreDataPort.scala 24:76:@46241.4]
  assign _T_45 = cnt > 5'h0; // @[StoreDataPort.scala 31:29:@46258.4]
  assign io_dataFromPrev_ready = cnt > 5'h0; // @[StoreDataPort.scala 32:25:@46262.4]
  assign io_storeDataEnable = _T_45 & io_dataFromPrev_valid; // @[StoreDataPort.scala 31:22:@46260.4]
  assign io_dataToStoreQueue = io_dataFromPrev_bits; // @[StoreDataPort.scala 30:23:@46257.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 5'h0;
    end else begin
      if (_T_30) begin
        cnt <= _T_33;
      end else begin
        if (_T_39) begin
          cnt <= _T_43;
        end
      end
    end
  end
endmodule
module LSQ_data( // @[:@46297.2]
  input         clock, // @[:@46298.4]
  input         reset, // @[:@46299.4]
  output [31:0] io_storeDataOut, // @[:@46300.4]
  output [31:0] io_storeAddrOut, // @[:@46300.4]
  output        io_storeEnable, // @[:@46300.4]
  input         io_memIsReadyForStores, // @[:@46300.4]
  input  [31:0] io_loadDataIn, // @[:@46300.4]
  output [31:0] io_loadAddrOut, // @[:@46300.4]
  output        io_loadEnable, // @[:@46300.4]
  input         io_memIsReadyForLoads, // @[:@46300.4]
  input         io_bbpValids_0, // @[:@46300.4]
  input         io_bbpValids_1, // @[:@46300.4]
  output        io_bbReadyToPrevs_0, // @[:@46300.4]
  output        io_bbReadyToPrevs_1, // @[:@46300.4]
  output        io_rdPortsPrev_0_ready, // @[:@46300.4]
  input         io_rdPortsPrev_0_valid, // @[:@46300.4]
  input  [31:0] io_rdPortsPrev_0_bits, // @[:@46300.4]
  output        io_rdPortsPrev_1_ready, // @[:@46300.4]
  input         io_rdPortsPrev_1_valid, // @[:@46300.4]
  input  [31:0] io_rdPortsPrev_1_bits, // @[:@46300.4]
  input         io_rdPortsNext_0_ready, // @[:@46300.4]
  output        io_rdPortsNext_0_valid, // @[:@46300.4]
  output [31:0] io_rdPortsNext_0_bits, // @[:@46300.4]
  input         io_rdPortsNext_1_ready, // @[:@46300.4]
  output        io_rdPortsNext_1_valid, // @[:@46300.4]
  output [31:0] io_rdPortsNext_1_bits, // @[:@46300.4]
  output        io_wrAddrPorts_0_ready, // @[:@46300.4]
  input         io_wrAddrPorts_0_valid, // @[:@46300.4]
  input  [31:0] io_wrAddrPorts_0_bits, // @[:@46300.4]
  output        io_wrDataPorts_0_ready, // @[:@46300.4]
  input         io_wrDataPorts_0_valid, // @[:@46300.4]
  input  [31:0] io_wrDataPorts_0_bits, // @[:@46300.4]
  output        io_Empty_Valid // @[:@46300.4]
);
  wire  storeQ_clock; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_reset; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_bbStart; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_bbStoreOffsets_0; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_bbStoreOffsets_1; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_bbStoreOffsets_2; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_bbStoreOffsets_3; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_bbStoreOffsets_4; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_bbStoreOffsets_5; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_bbStoreOffsets_6; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_bbStoreOffsets_7; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_bbStoreOffsets_8; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_bbStoreOffsets_9; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_bbStoreOffsets_10; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_bbStoreOffsets_11; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_bbStoreOffsets_12; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_bbStoreOffsets_13; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_bbStoreOffsets_14; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_bbStoreOffsets_15; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [1:0] storeQ_io_bbNumStores; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_storeTail; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_storeHead; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeEmpty; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_loadTail; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [3:0] storeQ_io_loadHead; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadEmpty; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadAddressDone_0; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadAddressDone_1; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadAddressDone_2; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadAddressDone_3; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadAddressDone_4; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadAddressDone_5; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadAddressDone_6; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadAddressDone_7; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadAddressDone_8; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadAddressDone_9; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadAddressDone_10; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadAddressDone_11; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadAddressDone_12; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadAddressDone_13; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadAddressDone_14; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadAddressDone_15; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadDataDone_0; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadDataDone_1; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadDataDone_2; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadDataDone_3; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadDataDone_4; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadDataDone_5; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadDataDone_6; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadDataDone_7; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadDataDone_8; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadDataDone_9; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadDataDone_10; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadDataDone_11; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadDataDone_12; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadDataDone_13; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadDataDone_14; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_loadDataDone_15; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_loadAddressQueue_0; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_loadAddressQueue_1; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_loadAddressQueue_2; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_loadAddressQueue_3; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_loadAddressQueue_4; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_loadAddressQueue_5; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_loadAddressQueue_6; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_loadAddressQueue_7; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_loadAddressQueue_8; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_loadAddressQueue_9; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_loadAddressQueue_10; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_loadAddressQueue_11; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_loadAddressQueue_12; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_loadAddressQueue_13; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_loadAddressQueue_14; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_loadAddressQueue_15; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeAddrDone_0; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeAddrDone_1; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeAddrDone_2; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeAddrDone_3; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeAddrDone_4; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeAddrDone_5; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeAddrDone_6; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeAddrDone_7; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeAddrDone_8; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeAddrDone_9; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeAddrDone_10; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeAddrDone_11; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeAddrDone_12; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeAddrDone_13; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeAddrDone_14; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeAddrDone_15; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeDataDone_0; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeDataDone_1; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeDataDone_2; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeDataDone_3; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeDataDone_4; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeDataDone_5; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeDataDone_6; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeDataDone_7; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeDataDone_8; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeDataDone_9; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeDataDone_10; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeDataDone_11; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeDataDone_12; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeDataDone_13; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeDataDone_14; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeDataDone_15; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeAddrQueue_0; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeAddrQueue_1; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeAddrQueue_2; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeAddrQueue_3; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeAddrQueue_4; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeAddrQueue_5; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeAddrQueue_6; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeAddrQueue_7; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeAddrQueue_8; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeAddrQueue_9; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeAddrQueue_10; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeAddrQueue_11; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeAddrQueue_12; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeAddrQueue_13; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeAddrQueue_14; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeAddrQueue_15; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeDataQueue_0; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeDataQueue_1; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeDataQueue_2; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeDataQueue_3; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeDataQueue_4; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeDataQueue_5; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeDataQueue_6; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeDataQueue_7; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeDataQueue_8; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeDataQueue_9; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeDataQueue_10; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeDataQueue_11; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeDataQueue_12; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeDataQueue_13; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeDataQueue_14; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeDataQueue_15; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeDataEnable_0; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_dataFromStorePorts_0; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeAddrEnable_0; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_addressFromStorePorts_0; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeAddrToMem; // @[LSQBRAM.scala 72:22:@46331.4]
  wire [31:0] storeQ_io_storeDataToMem; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_storeEnableToMem; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  storeQ_io_memIsReadyForStores; // @[LSQBRAM.scala 72:22:@46331.4]
  wire  loadQ_clock; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_reset; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_bbStart; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_bbLoadOffsets_0; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_bbLoadOffsets_1; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_bbLoadOffsets_2; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_bbLoadOffsets_3; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_bbLoadOffsets_4; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_bbLoadOffsets_5; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_bbLoadOffsets_6; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_bbLoadOffsets_7; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_bbLoadOffsets_8; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_bbLoadOffsets_9; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_bbLoadOffsets_10; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_bbLoadOffsets_11; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_bbLoadOffsets_12; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_bbLoadOffsets_13; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_bbLoadOffsets_14; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_bbLoadOffsets_15; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_bbLoadPorts_1; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [1:0] loadQ_io_bbNumLoads; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_loadTail; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_loadHead; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadEmpty; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_storeTail; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] loadQ_io_storeHead; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeEmpty; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeAddrDone_0; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeAddrDone_1; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeAddrDone_2; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeAddrDone_3; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeAddrDone_4; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeAddrDone_5; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeAddrDone_6; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeAddrDone_7; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeAddrDone_8; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeAddrDone_9; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeAddrDone_10; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeAddrDone_11; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeAddrDone_12; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeAddrDone_13; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeAddrDone_14; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeAddrDone_15; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeDataDone_0; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeDataDone_1; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeDataDone_2; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeDataDone_3; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeDataDone_4; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeDataDone_5; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeDataDone_6; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeDataDone_7; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeDataDone_8; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeDataDone_9; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeDataDone_10; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeDataDone_11; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeDataDone_12; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeDataDone_13; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeDataDone_14; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_storeDataDone_15; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeAddrQueue_0; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeAddrQueue_1; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeAddrQueue_2; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeAddrQueue_3; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeAddrQueue_4; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeAddrQueue_5; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeAddrQueue_6; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeAddrQueue_7; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeAddrQueue_8; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeAddrQueue_9; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeAddrQueue_10; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeAddrQueue_11; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeAddrQueue_12; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeAddrQueue_13; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeAddrQueue_14; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeAddrQueue_15; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeDataQueue_0; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeDataQueue_1; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeDataQueue_2; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeDataQueue_3; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeDataQueue_4; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeDataQueue_5; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeDataQueue_6; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeDataQueue_7; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeDataQueue_8; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeDataQueue_9; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeDataQueue_10; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeDataQueue_11; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeDataQueue_12; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeDataQueue_13; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeDataQueue_14; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_storeDataQueue_15; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrDone_0; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrDone_1; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrDone_2; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrDone_3; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrDone_4; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrDone_5; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrDone_6; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrDone_7; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrDone_8; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrDone_9; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrDone_10; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrDone_11; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrDone_12; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrDone_13; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrDone_14; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrDone_15; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadDataDone_0; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadDataDone_1; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadDataDone_2; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadDataDone_3; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadDataDone_4; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadDataDone_5; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadDataDone_6; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadDataDone_7; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadDataDone_8; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadDataDone_9; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadDataDone_10; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadDataDone_11; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadDataDone_12; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadDataDone_13; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadDataDone_14; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadDataDone_15; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadAddrQueue_0; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadAddrQueue_1; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadAddrQueue_2; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadAddrQueue_3; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadAddrQueue_4; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadAddrQueue_5; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadAddrQueue_6; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadAddrQueue_7; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadAddrQueue_8; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadAddrQueue_9; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadAddrQueue_10; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadAddrQueue_11; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadAddrQueue_12; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadAddrQueue_13; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadAddrQueue_14; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadAddrQueue_15; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrEnable_0; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadAddrEnable_1; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_addrFromLoadPorts_0; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_addrFromLoadPorts_1; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadPorts_0_ready; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadPorts_0_valid; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadPorts_0_bits; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadPorts_1_ready; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadPorts_1_valid; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadPorts_1_bits; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadDataFromMem; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [31:0] loadQ_io_loadAddrToMem; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_loadEnableToMem; // @[LSQBRAM.scala 73:21:@46334.4]
  wire  loadQ_io_memIsReadyForLoads; // @[LSQBRAM.scala 73:21:@46334.4]
  wire [3:0] GA_io_bbLoadOffsets_0; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbLoadOffsets_1; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbLoadOffsets_2; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbLoadOffsets_3; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbLoadOffsets_4; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbLoadOffsets_5; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbLoadOffsets_6; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbLoadOffsets_7; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbLoadOffsets_8; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbLoadOffsets_9; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbLoadOffsets_10; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbLoadOffsets_11; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbLoadOffsets_12; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbLoadOffsets_13; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbLoadOffsets_14; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbLoadOffsets_15; // @[LSQBRAM.scala 74:18:@46337.4]
  wire  GA_io_bbLoadPorts_1; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [1:0] GA_io_bbNumLoads; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_loadTail; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_loadHead; // @[LSQBRAM.scala 74:18:@46337.4]
  wire  GA_io_loadEmpty; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbStoreOffsets_0; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbStoreOffsets_1; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbStoreOffsets_2; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbStoreOffsets_3; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbStoreOffsets_4; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbStoreOffsets_5; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbStoreOffsets_6; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbStoreOffsets_7; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbStoreOffsets_8; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbStoreOffsets_9; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbStoreOffsets_10; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbStoreOffsets_11; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbStoreOffsets_12; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbStoreOffsets_13; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbStoreOffsets_14; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_bbStoreOffsets_15; // @[LSQBRAM.scala 74:18:@46337.4]
  wire  GA_io_bbNumStores; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_storeTail; // @[LSQBRAM.scala 74:18:@46337.4]
  wire [3:0] GA_io_storeHead; // @[LSQBRAM.scala 74:18:@46337.4]
  wire  GA_io_storeEmpty; // @[LSQBRAM.scala 74:18:@46337.4]
  wire  GA_io_bbStart; // @[LSQBRAM.scala 74:18:@46337.4]
  wire  GA_io_bbStartSignals_0; // @[LSQBRAM.scala 74:18:@46337.4]
  wire  GA_io_bbStartSignals_1; // @[LSQBRAM.scala 74:18:@46337.4]
  wire  GA_io_readyToPrevious_0; // @[LSQBRAM.scala 74:18:@46337.4]
  wire  GA_io_readyToPrevious_1; // @[LSQBRAM.scala 74:18:@46337.4]
  wire  GA_io_loadPortsEnable_0; // @[LSQBRAM.scala 74:18:@46337.4]
  wire  GA_io_loadPortsEnable_1; // @[LSQBRAM.scala 74:18:@46337.4]
  wire  GA_io_storePortsEnable_0; // @[LSQBRAM.scala 74:18:@46337.4]
  wire  LOAD_PORT_LSQ_data_clock; // @[LSQBRAM.scala 77:11:@46340.4]
  wire  LOAD_PORT_LSQ_data_reset; // @[LSQBRAM.scala 77:11:@46340.4]
  wire  LOAD_PORT_LSQ_data_io_addrFromPrev_ready; // @[LSQBRAM.scala 77:11:@46340.4]
  wire  LOAD_PORT_LSQ_data_io_addrFromPrev_valid; // @[LSQBRAM.scala 77:11:@46340.4]
  wire [31:0] LOAD_PORT_LSQ_data_io_addrFromPrev_bits; // @[LSQBRAM.scala 77:11:@46340.4]
  wire  LOAD_PORT_LSQ_data_io_portEnable; // @[LSQBRAM.scala 77:11:@46340.4]
  wire  LOAD_PORT_LSQ_data_io_dataToNext_ready; // @[LSQBRAM.scala 77:11:@46340.4]
  wire  LOAD_PORT_LSQ_data_io_dataToNext_valid; // @[LSQBRAM.scala 77:11:@46340.4]
  wire [31:0] LOAD_PORT_LSQ_data_io_dataToNext_bits; // @[LSQBRAM.scala 77:11:@46340.4]
  wire  LOAD_PORT_LSQ_data_io_loadAddrEnable; // @[LSQBRAM.scala 77:11:@46340.4]
  wire [31:0] LOAD_PORT_LSQ_data_io_addrToLoadQueue; // @[LSQBRAM.scala 77:11:@46340.4]
  wire  LOAD_PORT_LSQ_data_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 77:11:@46340.4]
  wire  LOAD_PORT_LSQ_data_io_dataFromLoadQueue_valid; // @[LSQBRAM.scala 77:11:@46340.4]
  wire [31:0] LOAD_PORT_LSQ_data_io_dataFromLoadQueue_bits; // @[LSQBRAM.scala 77:11:@46340.4]
  wire  LOAD_PORT_LSQ_data_1_clock; // @[LSQBRAM.scala 77:11:@46343.4]
  wire  LOAD_PORT_LSQ_data_1_reset; // @[LSQBRAM.scala 77:11:@46343.4]
  wire  LOAD_PORT_LSQ_data_1_io_addrFromPrev_ready; // @[LSQBRAM.scala 77:11:@46343.4]
  wire  LOAD_PORT_LSQ_data_1_io_addrFromPrev_valid; // @[LSQBRAM.scala 77:11:@46343.4]
  wire [31:0] LOAD_PORT_LSQ_data_1_io_addrFromPrev_bits; // @[LSQBRAM.scala 77:11:@46343.4]
  wire  LOAD_PORT_LSQ_data_1_io_portEnable; // @[LSQBRAM.scala 77:11:@46343.4]
  wire  LOAD_PORT_LSQ_data_1_io_dataToNext_ready; // @[LSQBRAM.scala 77:11:@46343.4]
  wire  LOAD_PORT_LSQ_data_1_io_dataToNext_valid; // @[LSQBRAM.scala 77:11:@46343.4]
  wire [31:0] LOAD_PORT_LSQ_data_1_io_dataToNext_bits; // @[LSQBRAM.scala 77:11:@46343.4]
  wire  LOAD_PORT_LSQ_data_1_io_loadAddrEnable; // @[LSQBRAM.scala 77:11:@46343.4]
  wire [31:0] LOAD_PORT_LSQ_data_1_io_addrToLoadQueue; // @[LSQBRAM.scala 77:11:@46343.4]
  wire  LOAD_PORT_LSQ_data_1_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 77:11:@46343.4]
  wire  LOAD_PORT_LSQ_data_1_io_dataFromLoadQueue_valid; // @[LSQBRAM.scala 77:11:@46343.4]
  wire [31:0] LOAD_PORT_LSQ_data_1_io_dataFromLoadQueue_bits; // @[LSQBRAM.scala 77:11:@46343.4]
  wire  STORE_DATA_PORT_LSQ_data_clock; // @[LSQBRAM.scala 80:11:@46371.4]
  wire  STORE_DATA_PORT_LSQ_data_reset; // @[LSQBRAM.scala 80:11:@46371.4]
  wire  STORE_DATA_PORT_LSQ_data_io_dataFromPrev_ready; // @[LSQBRAM.scala 80:11:@46371.4]
  wire  STORE_DATA_PORT_LSQ_data_io_dataFromPrev_valid; // @[LSQBRAM.scala 80:11:@46371.4]
  wire [31:0] STORE_DATA_PORT_LSQ_data_io_dataFromPrev_bits; // @[LSQBRAM.scala 80:11:@46371.4]
  wire  STORE_DATA_PORT_LSQ_data_io_portEnable; // @[LSQBRAM.scala 80:11:@46371.4]
  wire  STORE_DATA_PORT_LSQ_data_io_storeDataEnable; // @[LSQBRAM.scala 80:11:@46371.4]
  wire [31:0] STORE_DATA_PORT_LSQ_data_io_dataToStoreQueue; // @[LSQBRAM.scala 80:11:@46371.4]
  wire  STORE_ADDR_PORT_LSQ_data_clock; // @[LSQBRAM.scala 83:11:@46381.4]
  wire  STORE_ADDR_PORT_LSQ_data_reset; // @[LSQBRAM.scala 83:11:@46381.4]
  wire  STORE_ADDR_PORT_LSQ_data_io_dataFromPrev_ready; // @[LSQBRAM.scala 83:11:@46381.4]
  wire  STORE_ADDR_PORT_LSQ_data_io_dataFromPrev_valid; // @[LSQBRAM.scala 83:11:@46381.4]
  wire [31:0] STORE_ADDR_PORT_LSQ_data_io_dataFromPrev_bits; // @[LSQBRAM.scala 83:11:@46381.4]
  wire  STORE_ADDR_PORT_LSQ_data_io_portEnable; // @[LSQBRAM.scala 83:11:@46381.4]
  wire  STORE_ADDR_PORT_LSQ_data_io_storeDataEnable; // @[LSQBRAM.scala 83:11:@46381.4]
  wire [31:0] STORE_ADDR_PORT_LSQ_data_io_dataToStoreQueue; // @[LSQBRAM.scala 83:11:@46381.4]
  wire  storeEmpty; // @[LSQBRAM.scala 46:24:@46307.4 LSQBRAM.scala 151:14:@46726.4]
  wire  loadEmpty; // @[LSQBRAM.scala 52:23:@46313.4 LSQBRAM.scala 119:13:@46576.4]
  wire [15:0] storeTail; // @[LSQBRAM.scala 44:23:@46305.4 LSQBRAM.scala 149:13:@46724.4]
  wire [15:0] storeHead; // @[LSQBRAM.scala 45:23:@46306.4 LSQBRAM.scala 150:13:@46725.4]
  wire [15:0] loadTail; // @[LSQBRAM.scala 50:22:@46311.4 LSQBRAM.scala 117:12:@46574.4]
  wire [15:0] loadHead; // @[LSQBRAM.scala 51:22:@46312.4 LSQBRAM.scala 118:12:@46575.4]
  STORE_QUEUE_LSQ_data storeQ ( // @[LSQBRAM.scala 72:22:@46331.4]
    .clock(storeQ_clock),
    .reset(storeQ_reset),
    .io_bbStart(storeQ_io_bbStart),
    .io_bbStoreOffsets_0(storeQ_io_bbStoreOffsets_0),
    .io_bbStoreOffsets_1(storeQ_io_bbStoreOffsets_1),
    .io_bbStoreOffsets_2(storeQ_io_bbStoreOffsets_2),
    .io_bbStoreOffsets_3(storeQ_io_bbStoreOffsets_3),
    .io_bbStoreOffsets_4(storeQ_io_bbStoreOffsets_4),
    .io_bbStoreOffsets_5(storeQ_io_bbStoreOffsets_5),
    .io_bbStoreOffsets_6(storeQ_io_bbStoreOffsets_6),
    .io_bbStoreOffsets_7(storeQ_io_bbStoreOffsets_7),
    .io_bbStoreOffsets_8(storeQ_io_bbStoreOffsets_8),
    .io_bbStoreOffsets_9(storeQ_io_bbStoreOffsets_9),
    .io_bbStoreOffsets_10(storeQ_io_bbStoreOffsets_10),
    .io_bbStoreOffsets_11(storeQ_io_bbStoreOffsets_11),
    .io_bbStoreOffsets_12(storeQ_io_bbStoreOffsets_12),
    .io_bbStoreOffsets_13(storeQ_io_bbStoreOffsets_13),
    .io_bbStoreOffsets_14(storeQ_io_bbStoreOffsets_14),
    .io_bbStoreOffsets_15(storeQ_io_bbStoreOffsets_15),
    .io_bbNumStores(storeQ_io_bbNumStores),
    .io_storeTail(storeQ_io_storeTail),
    .io_storeHead(storeQ_io_storeHead),
    .io_storeEmpty(storeQ_io_storeEmpty),
    .io_loadTail(storeQ_io_loadTail),
    .io_loadHead(storeQ_io_loadHead),
    .io_loadEmpty(storeQ_io_loadEmpty),
    .io_loadAddressDone_0(storeQ_io_loadAddressDone_0),
    .io_loadAddressDone_1(storeQ_io_loadAddressDone_1),
    .io_loadAddressDone_2(storeQ_io_loadAddressDone_2),
    .io_loadAddressDone_3(storeQ_io_loadAddressDone_3),
    .io_loadAddressDone_4(storeQ_io_loadAddressDone_4),
    .io_loadAddressDone_5(storeQ_io_loadAddressDone_5),
    .io_loadAddressDone_6(storeQ_io_loadAddressDone_6),
    .io_loadAddressDone_7(storeQ_io_loadAddressDone_7),
    .io_loadAddressDone_8(storeQ_io_loadAddressDone_8),
    .io_loadAddressDone_9(storeQ_io_loadAddressDone_9),
    .io_loadAddressDone_10(storeQ_io_loadAddressDone_10),
    .io_loadAddressDone_11(storeQ_io_loadAddressDone_11),
    .io_loadAddressDone_12(storeQ_io_loadAddressDone_12),
    .io_loadAddressDone_13(storeQ_io_loadAddressDone_13),
    .io_loadAddressDone_14(storeQ_io_loadAddressDone_14),
    .io_loadAddressDone_15(storeQ_io_loadAddressDone_15),
    .io_loadDataDone_0(storeQ_io_loadDataDone_0),
    .io_loadDataDone_1(storeQ_io_loadDataDone_1),
    .io_loadDataDone_2(storeQ_io_loadDataDone_2),
    .io_loadDataDone_3(storeQ_io_loadDataDone_3),
    .io_loadDataDone_4(storeQ_io_loadDataDone_4),
    .io_loadDataDone_5(storeQ_io_loadDataDone_5),
    .io_loadDataDone_6(storeQ_io_loadDataDone_6),
    .io_loadDataDone_7(storeQ_io_loadDataDone_7),
    .io_loadDataDone_8(storeQ_io_loadDataDone_8),
    .io_loadDataDone_9(storeQ_io_loadDataDone_9),
    .io_loadDataDone_10(storeQ_io_loadDataDone_10),
    .io_loadDataDone_11(storeQ_io_loadDataDone_11),
    .io_loadDataDone_12(storeQ_io_loadDataDone_12),
    .io_loadDataDone_13(storeQ_io_loadDataDone_13),
    .io_loadDataDone_14(storeQ_io_loadDataDone_14),
    .io_loadDataDone_15(storeQ_io_loadDataDone_15),
    .io_loadAddressQueue_0(storeQ_io_loadAddressQueue_0),
    .io_loadAddressQueue_1(storeQ_io_loadAddressQueue_1),
    .io_loadAddressQueue_2(storeQ_io_loadAddressQueue_2),
    .io_loadAddressQueue_3(storeQ_io_loadAddressQueue_3),
    .io_loadAddressQueue_4(storeQ_io_loadAddressQueue_4),
    .io_loadAddressQueue_5(storeQ_io_loadAddressQueue_5),
    .io_loadAddressQueue_6(storeQ_io_loadAddressQueue_6),
    .io_loadAddressQueue_7(storeQ_io_loadAddressQueue_7),
    .io_loadAddressQueue_8(storeQ_io_loadAddressQueue_8),
    .io_loadAddressQueue_9(storeQ_io_loadAddressQueue_9),
    .io_loadAddressQueue_10(storeQ_io_loadAddressQueue_10),
    .io_loadAddressQueue_11(storeQ_io_loadAddressQueue_11),
    .io_loadAddressQueue_12(storeQ_io_loadAddressQueue_12),
    .io_loadAddressQueue_13(storeQ_io_loadAddressQueue_13),
    .io_loadAddressQueue_14(storeQ_io_loadAddressQueue_14),
    .io_loadAddressQueue_15(storeQ_io_loadAddressQueue_15),
    .io_storeAddrDone_0(storeQ_io_storeAddrDone_0),
    .io_storeAddrDone_1(storeQ_io_storeAddrDone_1),
    .io_storeAddrDone_2(storeQ_io_storeAddrDone_2),
    .io_storeAddrDone_3(storeQ_io_storeAddrDone_3),
    .io_storeAddrDone_4(storeQ_io_storeAddrDone_4),
    .io_storeAddrDone_5(storeQ_io_storeAddrDone_5),
    .io_storeAddrDone_6(storeQ_io_storeAddrDone_6),
    .io_storeAddrDone_7(storeQ_io_storeAddrDone_7),
    .io_storeAddrDone_8(storeQ_io_storeAddrDone_8),
    .io_storeAddrDone_9(storeQ_io_storeAddrDone_9),
    .io_storeAddrDone_10(storeQ_io_storeAddrDone_10),
    .io_storeAddrDone_11(storeQ_io_storeAddrDone_11),
    .io_storeAddrDone_12(storeQ_io_storeAddrDone_12),
    .io_storeAddrDone_13(storeQ_io_storeAddrDone_13),
    .io_storeAddrDone_14(storeQ_io_storeAddrDone_14),
    .io_storeAddrDone_15(storeQ_io_storeAddrDone_15),
    .io_storeDataDone_0(storeQ_io_storeDataDone_0),
    .io_storeDataDone_1(storeQ_io_storeDataDone_1),
    .io_storeDataDone_2(storeQ_io_storeDataDone_2),
    .io_storeDataDone_3(storeQ_io_storeDataDone_3),
    .io_storeDataDone_4(storeQ_io_storeDataDone_4),
    .io_storeDataDone_5(storeQ_io_storeDataDone_5),
    .io_storeDataDone_6(storeQ_io_storeDataDone_6),
    .io_storeDataDone_7(storeQ_io_storeDataDone_7),
    .io_storeDataDone_8(storeQ_io_storeDataDone_8),
    .io_storeDataDone_9(storeQ_io_storeDataDone_9),
    .io_storeDataDone_10(storeQ_io_storeDataDone_10),
    .io_storeDataDone_11(storeQ_io_storeDataDone_11),
    .io_storeDataDone_12(storeQ_io_storeDataDone_12),
    .io_storeDataDone_13(storeQ_io_storeDataDone_13),
    .io_storeDataDone_14(storeQ_io_storeDataDone_14),
    .io_storeDataDone_15(storeQ_io_storeDataDone_15),
    .io_storeAddrQueue_0(storeQ_io_storeAddrQueue_0),
    .io_storeAddrQueue_1(storeQ_io_storeAddrQueue_1),
    .io_storeAddrQueue_2(storeQ_io_storeAddrQueue_2),
    .io_storeAddrQueue_3(storeQ_io_storeAddrQueue_3),
    .io_storeAddrQueue_4(storeQ_io_storeAddrQueue_4),
    .io_storeAddrQueue_5(storeQ_io_storeAddrQueue_5),
    .io_storeAddrQueue_6(storeQ_io_storeAddrQueue_6),
    .io_storeAddrQueue_7(storeQ_io_storeAddrQueue_7),
    .io_storeAddrQueue_8(storeQ_io_storeAddrQueue_8),
    .io_storeAddrQueue_9(storeQ_io_storeAddrQueue_9),
    .io_storeAddrQueue_10(storeQ_io_storeAddrQueue_10),
    .io_storeAddrQueue_11(storeQ_io_storeAddrQueue_11),
    .io_storeAddrQueue_12(storeQ_io_storeAddrQueue_12),
    .io_storeAddrQueue_13(storeQ_io_storeAddrQueue_13),
    .io_storeAddrQueue_14(storeQ_io_storeAddrQueue_14),
    .io_storeAddrQueue_15(storeQ_io_storeAddrQueue_15),
    .io_storeDataQueue_0(storeQ_io_storeDataQueue_0),
    .io_storeDataQueue_1(storeQ_io_storeDataQueue_1),
    .io_storeDataQueue_2(storeQ_io_storeDataQueue_2),
    .io_storeDataQueue_3(storeQ_io_storeDataQueue_3),
    .io_storeDataQueue_4(storeQ_io_storeDataQueue_4),
    .io_storeDataQueue_5(storeQ_io_storeDataQueue_5),
    .io_storeDataQueue_6(storeQ_io_storeDataQueue_6),
    .io_storeDataQueue_7(storeQ_io_storeDataQueue_7),
    .io_storeDataQueue_8(storeQ_io_storeDataQueue_8),
    .io_storeDataQueue_9(storeQ_io_storeDataQueue_9),
    .io_storeDataQueue_10(storeQ_io_storeDataQueue_10),
    .io_storeDataQueue_11(storeQ_io_storeDataQueue_11),
    .io_storeDataQueue_12(storeQ_io_storeDataQueue_12),
    .io_storeDataQueue_13(storeQ_io_storeDataQueue_13),
    .io_storeDataQueue_14(storeQ_io_storeDataQueue_14),
    .io_storeDataQueue_15(storeQ_io_storeDataQueue_15),
    .io_storeDataEnable_0(storeQ_io_storeDataEnable_0),
    .io_dataFromStorePorts_0(storeQ_io_dataFromStorePorts_0),
    .io_storeAddrEnable_0(storeQ_io_storeAddrEnable_0),
    .io_addressFromStorePorts_0(storeQ_io_addressFromStorePorts_0),
    .io_storeAddrToMem(storeQ_io_storeAddrToMem),
    .io_storeDataToMem(storeQ_io_storeDataToMem),
    .io_storeEnableToMem(storeQ_io_storeEnableToMem),
    .io_memIsReadyForStores(storeQ_io_memIsReadyForStores)
  );
  LOAD_QUEUE_LSQ_data loadQ ( // @[LSQBRAM.scala 73:21:@46334.4]
    .clock(loadQ_clock),
    .reset(loadQ_reset),
    .io_bbStart(loadQ_io_bbStart),
    .io_bbLoadOffsets_0(loadQ_io_bbLoadOffsets_0),
    .io_bbLoadOffsets_1(loadQ_io_bbLoadOffsets_1),
    .io_bbLoadOffsets_2(loadQ_io_bbLoadOffsets_2),
    .io_bbLoadOffsets_3(loadQ_io_bbLoadOffsets_3),
    .io_bbLoadOffsets_4(loadQ_io_bbLoadOffsets_4),
    .io_bbLoadOffsets_5(loadQ_io_bbLoadOffsets_5),
    .io_bbLoadOffsets_6(loadQ_io_bbLoadOffsets_6),
    .io_bbLoadOffsets_7(loadQ_io_bbLoadOffsets_7),
    .io_bbLoadOffsets_8(loadQ_io_bbLoadOffsets_8),
    .io_bbLoadOffsets_9(loadQ_io_bbLoadOffsets_9),
    .io_bbLoadOffsets_10(loadQ_io_bbLoadOffsets_10),
    .io_bbLoadOffsets_11(loadQ_io_bbLoadOffsets_11),
    .io_bbLoadOffsets_12(loadQ_io_bbLoadOffsets_12),
    .io_bbLoadOffsets_13(loadQ_io_bbLoadOffsets_13),
    .io_bbLoadOffsets_14(loadQ_io_bbLoadOffsets_14),
    .io_bbLoadOffsets_15(loadQ_io_bbLoadOffsets_15),
    .io_bbLoadPorts_1(loadQ_io_bbLoadPorts_1),
    .io_bbNumLoads(loadQ_io_bbNumLoads),
    .io_loadTail(loadQ_io_loadTail),
    .io_loadHead(loadQ_io_loadHead),
    .io_loadEmpty(loadQ_io_loadEmpty),
    .io_storeTail(loadQ_io_storeTail),
    .io_storeHead(loadQ_io_storeHead),
    .io_storeEmpty(loadQ_io_storeEmpty),
    .io_storeAddrDone_0(loadQ_io_storeAddrDone_0),
    .io_storeAddrDone_1(loadQ_io_storeAddrDone_1),
    .io_storeAddrDone_2(loadQ_io_storeAddrDone_2),
    .io_storeAddrDone_3(loadQ_io_storeAddrDone_3),
    .io_storeAddrDone_4(loadQ_io_storeAddrDone_4),
    .io_storeAddrDone_5(loadQ_io_storeAddrDone_5),
    .io_storeAddrDone_6(loadQ_io_storeAddrDone_6),
    .io_storeAddrDone_7(loadQ_io_storeAddrDone_7),
    .io_storeAddrDone_8(loadQ_io_storeAddrDone_8),
    .io_storeAddrDone_9(loadQ_io_storeAddrDone_9),
    .io_storeAddrDone_10(loadQ_io_storeAddrDone_10),
    .io_storeAddrDone_11(loadQ_io_storeAddrDone_11),
    .io_storeAddrDone_12(loadQ_io_storeAddrDone_12),
    .io_storeAddrDone_13(loadQ_io_storeAddrDone_13),
    .io_storeAddrDone_14(loadQ_io_storeAddrDone_14),
    .io_storeAddrDone_15(loadQ_io_storeAddrDone_15),
    .io_storeDataDone_0(loadQ_io_storeDataDone_0),
    .io_storeDataDone_1(loadQ_io_storeDataDone_1),
    .io_storeDataDone_2(loadQ_io_storeDataDone_2),
    .io_storeDataDone_3(loadQ_io_storeDataDone_3),
    .io_storeDataDone_4(loadQ_io_storeDataDone_4),
    .io_storeDataDone_5(loadQ_io_storeDataDone_5),
    .io_storeDataDone_6(loadQ_io_storeDataDone_6),
    .io_storeDataDone_7(loadQ_io_storeDataDone_7),
    .io_storeDataDone_8(loadQ_io_storeDataDone_8),
    .io_storeDataDone_9(loadQ_io_storeDataDone_9),
    .io_storeDataDone_10(loadQ_io_storeDataDone_10),
    .io_storeDataDone_11(loadQ_io_storeDataDone_11),
    .io_storeDataDone_12(loadQ_io_storeDataDone_12),
    .io_storeDataDone_13(loadQ_io_storeDataDone_13),
    .io_storeDataDone_14(loadQ_io_storeDataDone_14),
    .io_storeDataDone_15(loadQ_io_storeDataDone_15),
    .io_storeAddrQueue_0(loadQ_io_storeAddrQueue_0),
    .io_storeAddrQueue_1(loadQ_io_storeAddrQueue_1),
    .io_storeAddrQueue_2(loadQ_io_storeAddrQueue_2),
    .io_storeAddrQueue_3(loadQ_io_storeAddrQueue_3),
    .io_storeAddrQueue_4(loadQ_io_storeAddrQueue_4),
    .io_storeAddrQueue_5(loadQ_io_storeAddrQueue_5),
    .io_storeAddrQueue_6(loadQ_io_storeAddrQueue_6),
    .io_storeAddrQueue_7(loadQ_io_storeAddrQueue_7),
    .io_storeAddrQueue_8(loadQ_io_storeAddrQueue_8),
    .io_storeAddrQueue_9(loadQ_io_storeAddrQueue_9),
    .io_storeAddrQueue_10(loadQ_io_storeAddrQueue_10),
    .io_storeAddrQueue_11(loadQ_io_storeAddrQueue_11),
    .io_storeAddrQueue_12(loadQ_io_storeAddrQueue_12),
    .io_storeAddrQueue_13(loadQ_io_storeAddrQueue_13),
    .io_storeAddrQueue_14(loadQ_io_storeAddrQueue_14),
    .io_storeAddrQueue_15(loadQ_io_storeAddrQueue_15),
    .io_storeDataQueue_0(loadQ_io_storeDataQueue_0),
    .io_storeDataQueue_1(loadQ_io_storeDataQueue_1),
    .io_storeDataQueue_2(loadQ_io_storeDataQueue_2),
    .io_storeDataQueue_3(loadQ_io_storeDataQueue_3),
    .io_storeDataQueue_4(loadQ_io_storeDataQueue_4),
    .io_storeDataQueue_5(loadQ_io_storeDataQueue_5),
    .io_storeDataQueue_6(loadQ_io_storeDataQueue_6),
    .io_storeDataQueue_7(loadQ_io_storeDataQueue_7),
    .io_storeDataQueue_8(loadQ_io_storeDataQueue_8),
    .io_storeDataQueue_9(loadQ_io_storeDataQueue_9),
    .io_storeDataQueue_10(loadQ_io_storeDataQueue_10),
    .io_storeDataQueue_11(loadQ_io_storeDataQueue_11),
    .io_storeDataQueue_12(loadQ_io_storeDataQueue_12),
    .io_storeDataQueue_13(loadQ_io_storeDataQueue_13),
    .io_storeDataQueue_14(loadQ_io_storeDataQueue_14),
    .io_storeDataQueue_15(loadQ_io_storeDataQueue_15),
    .io_loadAddrDone_0(loadQ_io_loadAddrDone_0),
    .io_loadAddrDone_1(loadQ_io_loadAddrDone_1),
    .io_loadAddrDone_2(loadQ_io_loadAddrDone_2),
    .io_loadAddrDone_3(loadQ_io_loadAddrDone_3),
    .io_loadAddrDone_4(loadQ_io_loadAddrDone_4),
    .io_loadAddrDone_5(loadQ_io_loadAddrDone_5),
    .io_loadAddrDone_6(loadQ_io_loadAddrDone_6),
    .io_loadAddrDone_7(loadQ_io_loadAddrDone_7),
    .io_loadAddrDone_8(loadQ_io_loadAddrDone_8),
    .io_loadAddrDone_9(loadQ_io_loadAddrDone_9),
    .io_loadAddrDone_10(loadQ_io_loadAddrDone_10),
    .io_loadAddrDone_11(loadQ_io_loadAddrDone_11),
    .io_loadAddrDone_12(loadQ_io_loadAddrDone_12),
    .io_loadAddrDone_13(loadQ_io_loadAddrDone_13),
    .io_loadAddrDone_14(loadQ_io_loadAddrDone_14),
    .io_loadAddrDone_15(loadQ_io_loadAddrDone_15),
    .io_loadDataDone_0(loadQ_io_loadDataDone_0),
    .io_loadDataDone_1(loadQ_io_loadDataDone_1),
    .io_loadDataDone_2(loadQ_io_loadDataDone_2),
    .io_loadDataDone_3(loadQ_io_loadDataDone_3),
    .io_loadDataDone_4(loadQ_io_loadDataDone_4),
    .io_loadDataDone_5(loadQ_io_loadDataDone_5),
    .io_loadDataDone_6(loadQ_io_loadDataDone_6),
    .io_loadDataDone_7(loadQ_io_loadDataDone_7),
    .io_loadDataDone_8(loadQ_io_loadDataDone_8),
    .io_loadDataDone_9(loadQ_io_loadDataDone_9),
    .io_loadDataDone_10(loadQ_io_loadDataDone_10),
    .io_loadDataDone_11(loadQ_io_loadDataDone_11),
    .io_loadDataDone_12(loadQ_io_loadDataDone_12),
    .io_loadDataDone_13(loadQ_io_loadDataDone_13),
    .io_loadDataDone_14(loadQ_io_loadDataDone_14),
    .io_loadDataDone_15(loadQ_io_loadDataDone_15),
    .io_loadAddrQueue_0(loadQ_io_loadAddrQueue_0),
    .io_loadAddrQueue_1(loadQ_io_loadAddrQueue_1),
    .io_loadAddrQueue_2(loadQ_io_loadAddrQueue_2),
    .io_loadAddrQueue_3(loadQ_io_loadAddrQueue_3),
    .io_loadAddrQueue_4(loadQ_io_loadAddrQueue_4),
    .io_loadAddrQueue_5(loadQ_io_loadAddrQueue_5),
    .io_loadAddrQueue_6(loadQ_io_loadAddrQueue_6),
    .io_loadAddrQueue_7(loadQ_io_loadAddrQueue_7),
    .io_loadAddrQueue_8(loadQ_io_loadAddrQueue_8),
    .io_loadAddrQueue_9(loadQ_io_loadAddrQueue_9),
    .io_loadAddrQueue_10(loadQ_io_loadAddrQueue_10),
    .io_loadAddrQueue_11(loadQ_io_loadAddrQueue_11),
    .io_loadAddrQueue_12(loadQ_io_loadAddrQueue_12),
    .io_loadAddrQueue_13(loadQ_io_loadAddrQueue_13),
    .io_loadAddrQueue_14(loadQ_io_loadAddrQueue_14),
    .io_loadAddrQueue_15(loadQ_io_loadAddrQueue_15),
    .io_loadAddrEnable_0(loadQ_io_loadAddrEnable_0),
    .io_loadAddrEnable_1(loadQ_io_loadAddrEnable_1),
    .io_addrFromLoadPorts_0(loadQ_io_addrFromLoadPorts_0),
    .io_addrFromLoadPorts_1(loadQ_io_addrFromLoadPorts_1),
    .io_loadPorts_0_ready(loadQ_io_loadPorts_0_ready),
    .io_loadPorts_0_valid(loadQ_io_loadPorts_0_valid),
    .io_loadPorts_0_bits(loadQ_io_loadPorts_0_bits),
    .io_loadPorts_1_ready(loadQ_io_loadPorts_1_ready),
    .io_loadPorts_1_valid(loadQ_io_loadPorts_1_valid),
    .io_loadPorts_1_bits(loadQ_io_loadPorts_1_bits),
    .io_loadDataFromMem(loadQ_io_loadDataFromMem),
    .io_loadAddrToMem(loadQ_io_loadAddrToMem),
    .io_loadEnableToMem(loadQ_io_loadEnableToMem),
    .io_memIsReadyForLoads(loadQ_io_memIsReadyForLoads)
  );
  GROUP_ALLOCATOR_LSQ_data GA ( // @[LSQBRAM.scala 74:18:@46337.4]
    .io_bbLoadOffsets_0(GA_io_bbLoadOffsets_0),
    .io_bbLoadOffsets_1(GA_io_bbLoadOffsets_1),
    .io_bbLoadOffsets_2(GA_io_bbLoadOffsets_2),
    .io_bbLoadOffsets_3(GA_io_bbLoadOffsets_3),
    .io_bbLoadOffsets_4(GA_io_bbLoadOffsets_4),
    .io_bbLoadOffsets_5(GA_io_bbLoadOffsets_5),
    .io_bbLoadOffsets_6(GA_io_bbLoadOffsets_6),
    .io_bbLoadOffsets_7(GA_io_bbLoadOffsets_7),
    .io_bbLoadOffsets_8(GA_io_bbLoadOffsets_8),
    .io_bbLoadOffsets_9(GA_io_bbLoadOffsets_9),
    .io_bbLoadOffsets_10(GA_io_bbLoadOffsets_10),
    .io_bbLoadOffsets_11(GA_io_bbLoadOffsets_11),
    .io_bbLoadOffsets_12(GA_io_bbLoadOffsets_12),
    .io_bbLoadOffsets_13(GA_io_bbLoadOffsets_13),
    .io_bbLoadOffsets_14(GA_io_bbLoadOffsets_14),
    .io_bbLoadOffsets_15(GA_io_bbLoadOffsets_15),
    .io_bbLoadPorts_1(GA_io_bbLoadPorts_1),
    .io_bbNumLoads(GA_io_bbNumLoads),
    .io_loadTail(GA_io_loadTail),
    .io_loadHead(GA_io_loadHead),
    .io_loadEmpty(GA_io_loadEmpty),
    .io_bbStoreOffsets_0(GA_io_bbStoreOffsets_0),
    .io_bbStoreOffsets_1(GA_io_bbStoreOffsets_1),
    .io_bbStoreOffsets_2(GA_io_bbStoreOffsets_2),
    .io_bbStoreOffsets_3(GA_io_bbStoreOffsets_3),
    .io_bbStoreOffsets_4(GA_io_bbStoreOffsets_4),
    .io_bbStoreOffsets_5(GA_io_bbStoreOffsets_5),
    .io_bbStoreOffsets_6(GA_io_bbStoreOffsets_6),
    .io_bbStoreOffsets_7(GA_io_bbStoreOffsets_7),
    .io_bbStoreOffsets_8(GA_io_bbStoreOffsets_8),
    .io_bbStoreOffsets_9(GA_io_bbStoreOffsets_9),
    .io_bbStoreOffsets_10(GA_io_bbStoreOffsets_10),
    .io_bbStoreOffsets_11(GA_io_bbStoreOffsets_11),
    .io_bbStoreOffsets_12(GA_io_bbStoreOffsets_12),
    .io_bbStoreOffsets_13(GA_io_bbStoreOffsets_13),
    .io_bbStoreOffsets_14(GA_io_bbStoreOffsets_14),
    .io_bbStoreOffsets_15(GA_io_bbStoreOffsets_15),
    .io_bbNumStores(GA_io_bbNumStores),
    .io_storeTail(GA_io_storeTail),
    .io_storeHead(GA_io_storeHead),
    .io_storeEmpty(GA_io_storeEmpty),
    .io_bbStart(GA_io_bbStart),
    .io_bbStartSignals_0(GA_io_bbStartSignals_0),
    .io_bbStartSignals_1(GA_io_bbStartSignals_1),
    .io_readyToPrevious_0(GA_io_readyToPrevious_0),
    .io_readyToPrevious_1(GA_io_readyToPrevious_1),
    .io_loadPortsEnable_0(GA_io_loadPortsEnable_0),
    .io_loadPortsEnable_1(GA_io_loadPortsEnable_1),
    .io_storePortsEnable_0(GA_io_storePortsEnable_0)
  );
  LOAD_PORT_LSQ_data LOAD_PORT_LSQ_data ( // @[LSQBRAM.scala 77:11:@46340.4]
    .clock(LOAD_PORT_LSQ_data_clock),
    .reset(LOAD_PORT_LSQ_data_reset),
    .io_addrFromPrev_ready(LOAD_PORT_LSQ_data_io_addrFromPrev_ready),
    .io_addrFromPrev_valid(LOAD_PORT_LSQ_data_io_addrFromPrev_valid),
    .io_addrFromPrev_bits(LOAD_PORT_LSQ_data_io_addrFromPrev_bits),
    .io_portEnable(LOAD_PORT_LSQ_data_io_portEnable),
    .io_dataToNext_ready(LOAD_PORT_LSQ_data_io_dataToNext_ready),
    .io_dataToNext_valid(LOAD_PORT_LSQ_data_io_dataToNext_valid),
    .io_dataToNext_bits(LOAD_PORT_LSQ_data_io_dataToNext_bits),
    .io_loadAddrEnable(LOAD_PORT_LSQ_data_io_loadAddrEnable),
    .io_addrToLoadQueue(LOAD_PORT_LSQ_data_io_addrToLoadQueue),
    .io_dataFromLoadQueue_ready(LOAD_PORT_LSQ_data_io_dataFromLoadQueue_ready),
    .io_dataFromLoadQueue_valid(LOAD_PORT_LSQ_data_io_dataFromLoadQueue_valid),
    .io_dataFromLoadQueue_bits(LOAD_PORT_LSQ_data_io_dataFromLoadQueue_bits)
  );
  LOAD_PORT_LSQ_data LOAD_PORT_LSQ_data_1 ( // @[LSQBRAM.scala 77:11:@46343.4]
    .clock(LOAD_PORT_LSQ_data_1_clock),
    .reset(LOAD_PORT_LSQ_data_1_reset),
    .io_addrFromPrev_ready(LOAD_PORT_LSQ_data_1_io_addrFromPrev_ready),
    .io_addrFromPrev_valid(LOAD_PORT_LSQ_data_1_io_addrFromPrev_valid),
    .io_addrFromPrev_bits(LOAD_PORT_LSQ_data_1_io_addrFromPrev_bits),
    .io_portEnable(LOAD_PORT_LSQ_data_1_io_portEnable),
    .io_dataToNext_ready(LOAD_PORT_LSQ_data_1_io_dataToNext_ready),
    .io_dataToNext_valid(LOAD_PORT_LSQ_data_1_io_dataToNext_valid),
    .io_dataToNext_bits(LOAD_PORT_LSQ_data_1_io_dataToNext_bits),
    .io_loadAddrEnable(LOAD_PORT_LSQ_data_1_io_loadAddrEnable),
    .io_addrToLoadQueue(LOAD_PORT_LSQ_data_1_io_addrToLoadQueue),
    .io_dataFromLoadQueue_ready(LOAD_PORT_LSQ_data_1_io_dataFromLoadQueue_ready),
    .io_dataFromLoadQueue_valid(LOAD_PORT_LSQ_data_1_io_dataFromLoadQueue_valid),
    .io_dataFromLoadQueue_bits(LOAD_PORT_LSQ_data_1_io_dataFromLoadQueue_bits)
  );
  STORE_DATA_PORT_LSQ_data STORE_DATA_PORT_LSQ_data ( // @[LSQBRAM.scala 80:11:@46371.4]
    .clock(STORE_DATA_PORT_LSQ_data_clock),
    .reset(STORE_DATA_PORT_LSQ_data_reset),
    .io_dataFromPrev_ready(STORE_DATA_PORT_LSQ_data_io_dataFromPrev_ready),
    .io_dataFromPrev_valid(STORE_DATA_PORT_LSQ_data_io_dataFromPrev_valid),
    .io_dataFromPrev_bits(STORE_DATA_PORT_LSQ_data_io_dataFromPrev_bits),
    .io_portEnable(STORE_DATA_PORT_LSQ_data_io_portEnable),
    .io_storeDataEnable(STORE_DATA_PORT_LSQ_data_io_storeDataEnable),
    .io_dataToStoreQueue(STORE_DATA_PORT_LSQ_data_io_dataToStoreQueue)
  );
  STORE_DATA_PORT_LSQ_data STORE_ADDR_PORT_LSQ_data ( // @[LSQBRAM.scala 83:11:@46381.4]
    .clock(STORE_ADDR_PORT_LSQ_data_clock),
    .reset(STORE_ADDR_PORT_LSQ_data_reset),
    .io_dataFromPrev_ready(STORE_ADDR_PORT_LSQ_data_io_dataFromPrev_ready),
    .io_dataFromPrev_valid(STORE_ADDR_PORT_LSQ_data_io_dataFromPrev_valid),
    .io_dataFromPrev_bits(STORE_ADDR_PORT_LSQ_data_io_dataFromPrev_bits),
    .io_portEnable(STORE_ADDR_PORT_LSQ_data_io_portEnable),
    .io_storeDataEnable(STORE_ADDR_PORT_LSQ_data_io_storeDataEnable),
    .io_dataToStoreQueue(STORE_ADDR_PORT_LSQ_data_io_dataToStoreQueue)
  );
  assign storeEmpty = storeQ_io_storeEmpty; // @[LSQBRAM.scala 46:24:@46307.4 LSQBRAM.scala 151:14:@46726.4]
  assign loadEmpty = loadQ_io_loadEmpty; // @[LSQBRAM.scala 52:23:@46313.4 LSQBRAM.scala 119:13:@46576.4]
  assign storeTail = {{12'd0}, storeQ_io_storeTail}; // @[LSQBRAM.scala 44:23:@46305.4 LSQBRAM.scala 149:13:@46724.4]
  assign storeHead = {{12'd0}, storeQ_io_storeHead}; // @[LSQBRAM.scala 45:23:@46306.4 LSQBRAM.scala 150:13:@46725.4]
  assign loadTail = {{12'd0}, loadQ_io_loadTail}; // @[LSQBRAM.scala 50:22:@46311.4 LSQBRAM.scala 117:12:@46574.4]
  assign loadHead = {{12'd0}, loadQ_io_loadHead}; // @[LSQBRAM.scala 51:22:@46312.4 LSQBRAM.scala 118:12:@46575.4]
  assign io_storeDataOut = storeQ_io_storeDataToMem; // @[LSQBRAM.scala 161:19:@46796.4]
  assign io_storeAddrOut = storeQ_io_storeAddrToMem; // @[LSQBRAM.scala 160:19:@46795.4]
  assign io_storeEnable = storeQ_io_storeEnableToMem; // @[LSQBRAM.scala 162:18:@46797.4]
  assign io_loadAddrOut = loadQ_io_loadAddrToMem; // @[LSQBRAM.scala 135:18:@46637.4]
  assign io_loadEnable = loadQ_io_loadEnableToMem; // @[LSQBRAM.scala 136:17:@46638.4]
  assign io_bbReadyToPrevs_0 = GA_io_readyToPrevious_0; // @[LSQBRAM.scala 102:21:@46468.4]
  assign io_bbReadyToPrevs_1 = GA_io_readyToPrevious_1; // @[LSQBRAM.scala 102:21:@46469.4]
  assign io_rdPortsPrev_0_ready = LOAD_PORT_LSQ_data_io_addrFromPrev_ready; // @[LSQBRAM.scala 166:31:@46801.4]
  assign io_rdPortsPrev_1_ready = LOAD_PORT_LSQ_data_1_io_addrFromPrev_ready; // @[LSQBRAM.scala 166:31:@46813.4]
  assign io_rdPortsNext_0_valid = LOAD_PORT_LSQ_data_io_dataToNext_valid; // @[LSQBRAM.scala 168:23:@46804.4]
  assign io_rdPortsNext_0_bits = LOAD_PORT_LSQ_data_io_dataToNext_bits; // @[LSQBRAM.scala 168:23:@46803.4]
  assign io_rdPortsNext_1_valid = LOAD_PORT_LSQ_data_1_io_dataToNext_valid; // @[LSQBRAM.scala 168:23:@46816.4]
  assign io_rdPortsNext_1_bits = LOAD_PORT_LSQ_data_1_io_dataToNext_bits; // @[LSQBRAM.scala 168:23:@46815.4]
  assign io_wrAddrPorts_0_ready = STORE_ADDR_PORT_LSQ_data_io_dataFromPrev_ready; // @[LSQBRAM.scala 182:39:@46831.4]
  assign io_wrDataPorts_0_ready = STORE_DATA_PORT_LSQ_data_io_dataFromPrev_ready; // @[LSQBRAM.scala 177:36:@46825.4]
  assign io_Empty_Valid = storeEmpty & loadEmpty; // @[LSQBRAM.scala 86:18:@46392.4]
  assign storeQ_clock = clock; // @[:@46332.4]
  assign storeQ_reset = reset; // @[:@46333.4]
  assign storeQ_io_bbStart = GA_io_bbStart; // @[LSQBRAM.scala 145:21:@46690.4]
  assign storeQ_io_bbStoreOffsets_0 = GA_io_bbStoreOffsets_0; // @[LSQBRAM.scala 146:28:@46691.4]
  assign storeQ_io_bbStoreOffsets_1 = GA_io_bbStoreOffsets_1; // @[LSQBRAM.scala 146:28:@46692.4]
  assign storeQ_io_bbStoreOffsets_2 = GA_io_bbStoreOffsets_2; // @[LSQBRAM.scala 146:28:@46693.4]
  assign storeQ_io_bbStoreOffsets_3 = GA_io_bbStoreOffsets_3; // @[LSQBRAM.scala 146:28:@46694.4]
  assign storeQ_io_bbStoreOffsets_4 = GA_io_bbStoreOffsets_4; // @[LSQBRAM.scala 146:28:@46695.4]
  assign storeQ_io_bbStoreOffsets_5 = GA_io_bbStoreOffsets_5; // @[LSQBRAM.scala 146:28:@46696.4]
  assign storeQ_io_bbStoreOffsets_6 = GA_io_bbStoreOffsets_6; // @[LSQBRAM.scala 146:28:@46697.4]
  assign storeQ_io_bbStoreOffsets_7 = GA_io_bbStoreOffsets_7; // @[LSQBRAM.scala 146:28:@46698.4]
  assign storeQ_io_bbStoreOffsets_8 = GA_io_bbStoreOffsets_8; // @[LSQBRAM.scala 146:28:@46699.4]
  assign storeQ_io_bbStoreOffsets_9 = GA_io_bbStoreOffsets_9; // @[LSQBRAM.scala 146:28:@46700.4]
  assign storeQ_io_bbStoreOffsets_10 = GA_io_bbStoreOffsets_10; // @[LSQBRAM.scala 146:28:@46701.4]
  assign storeQ_io_bbStoreOffsets_11 = GA_io_bbStoreOffsets_11; // @[LSQBRAM.scala 146:28:@46702.4]
  assign storeQ_io_bbStoreOffsets_12 = GA_io_bbStoreOffsets_12; // @[LSQBRAM.scala 146:28:@46703.4]
  assign storeQ_io_bbStoreOffsets_13 = GA_io_bbStoreOffsets_13; // @[LSQBRAM.scala 146:28:@46704.4]
  assign storeQ_io_bbStoreOffsets_14 = GA_io_bbStoreOffsets_14; // @[LSQBRAM.scala 146:28:@46705.4]
  assign storeQ_io_bbStoreOffsets_15 = GA_io_bbStoreOffsets_15; // @[LSQBRAM.scala 146:28:@46706.4]
  assign storeQ_io_bbNumStores = {{1'd0}, GA_io_bbNumStores}; // @[LSQBRAM.scala 148:25:@46723.4]
  assign storeQ_io_loadTail = loadTail[3:0]; // @[LSQBRAM.scala 139:22:@46639.4]
  assign storeQ_io_loadHead = loadHead[3:0]; // @[LSQBRAM.scala 140:22:@46640.4]
  assign storeQ_io_loadEmpty = loadQ_io_loadEmpty; // @[LSQBRAM.scala 141:23:@46641.4]
  assign storeQ_io_loadAddressDone_0 = loadQ_io_loadAddrDone_0; // @[LSQBRAM.scala 142:29:@46642.4]
  assign storeQ_io_loadAddressDone_1 = loadQ_io_loadAddrDone_1; // @[LSQBRAM.scala 142:29:@46643.4]
  assign storeQ_io_loadAddressDone_2 = loadQ_io_loadAddrDone_2; // @[LSQBRAM.scala 142:29:@46644.4]
  assign storeQ_io_loadAddressDone_3 = loadQ_io_loadAddrDone_3; // @[LSQBRAM.scala 142:29:@46645.4]
  assign storeQ_io_loadAddressDone_4 = loadQ_io_loadAddrDone_4; // @[LSQBRAM.scala 142:29:@46646.4]
  assign storeQ_io_loadAddressDone_5 = loadQ_io_loadAddrDone_5; // @[LSQBRAM.scala 142:29:@46647.4]
  assign storeQ_io_loadAddressDone_6 = loadQ_io_loadAddrDone_6; // @[LSQBRAM.scala 142:29:@46648.4]
  assign storeQ_io_loadAddressDone_7 = loadQ_io_loadAddrDone_7; // @[LSQBRAM.scala 142:29:@46649.4]
  assign storeQ_io_loadAddressDone_8 = loadQ_io_loadAddrDone_8; // @[LSQBRAM.scala 142:29:@46650.4]
  assign storeQ_io_loadAddressDone_9 = loadQ_io_loadAddrDone_9; // @[LSQBRAM.scala 142:29:@46651.4]
  assign storeQ_io_loadAddressDone_10 = loadQ_io_loadAddrDone_10; // @[LSQBRAM.scala 142:29:@46652.4]
  assign storeQ_io_loadAddressDone_11 = loadQ_io_loadAddrDone_11; // @[LSQBRAM.scala 142:29:@46653.4]
  assign storeQ_io_loadAddressDone_12 = loadQ_io_loadAddrDone_12; // @[LSQBRAM.scala 142:29:@46654.4]
  assign storeQ_io_loadAddressDone_13 = loadQ_io_loadAddrDone_13; // @[LSQBRAM.scala 142:29:@46655.4]
  assign storeQ_io_loadAddressDone_14 = loadQ_io_loadAddrDone_14; // @[LSQBRAM.scala 142:29:@46656.4]
  assign storeQ_io_loadAddressDone_15 = loadQ_io_loadAddrDone_15; // @[LSQBRAM.scala 142:29:@46657.4]
  assign storeQ_io_loadDataDone_0 = loadQ_io_loadDataDone_0; // @[LSQBRAM.scala 143:26:@46658.4]
  assign storeQ_io_loadDataDone_1 = loadQ_io_loadDataDone_1; // @[LSQBRAM.scala 143:26:@46659.4]
  assign storeQ_io_loadDataDone_2 = loadQ_io_loadDataDone_2; // @[LSQBRAM.scala 143:26:@46660.4]
  assign storeQ_io_loadDataDone_3 = loadQ_io_loadDataDone_3; // @[LSQBRAM.scala 143:26:@46661.4]
  assign storeQ_io_loadDataDone_4 = loadQ_io_loadDataDone_4; // @[LSQBRAM.scala 143:26:@46662.4]
  assign storeQ_io_loadDataDone_5 = loadQ_io_loadDataDone_5; // @[LSQBRAM.scala 143:26:@46663.4]
  assign storeQ_io_loadDataDone_6 = loadQ_io_loadDataDone_6; // @[LSQBRAM.scala 143:26:@46664.4]
  assign storeQ_io_loadDataDone_7 = loadQ_io_loadDataDone_7; // @[LSQBRAM.scala 143:26:@46665.4]
  assign storeQ_io_loadDataDone_8 = loadQ_io_loadDataDone_8; // @[LSQBRAM.scala 143:26:@46666.4]
  assign storeQ_io_loadDataDone_9 = loadQ_io_loadDataDone_9; // @[LSQBRAM.scala 143:26:@46667.4]
  assign storeQ_io_loadDataDone_10 = loadQ_io_loadDataDone_10; // @[LSQBRAM.scala 143:26:@46668.4]
  assign storeQ_io_loadDataDone_11 = loadQ_io_loadDataDone_11; // @[LSQBRAM.scala 143:26:@46669.4]
  assign storeQ_io_loadDataDone_12 = loadQ_io_loadDataDone_12; // @[LSQBRAM.scala 143:26:@46670.4]
  assign storeQ_io_loadDataDone_13 = loadQ_io_loadDataDone_13; // @[LSQBRAM.scala 143:26:@46671.4]
  assign storeQ_io_loadDataDone_14 = loadQ_io_loadDataDone_14; // @[LSQBRAM.scala 143:26:@46672.4]
  assign storeQ_io_loadDataDone_15 = loadQ_io_loadDataDone_15; // @[LSQBRAM.scala 143:26:@46673.4]
  assign storeQ_io_loadAddressQueue_0 = loadQ_io_loadAddrQueue_0; // @[LSQBRAM.scala 144:30:@46674.4]
  assign storeQ_io_loadAddressQueue_1 = loadQ_io_loadAddrQueue_1; // @[LSQBRAM.scala 144:30:@46675.4]
  assign storeQ_io_loadAddressQueue_2 = loadQ_io_loadAddrQueue_2; // @[LSQBRAM.scala 144:30:@46676.4]
  assign storeQ_io_loadAddressQueue_3 = loadQ_io_loadAddrQueue_3; // @[LSQBRAM.scala 144:30:@46677.4]
  assign storeQ_io_loadAddressQueue_4 = loadQ_io_loadAddrQueue_4; // @[LSQBRAM.scala 144:30:@46678.4]
  assign storeQ_io_loadAddressQueue_5 = loadQ_io_loadAddrQueue_5; // @[LSQBRAM.scala 144:30:@46679.4]
  assign storeQ_io_loadAddressQueue_6 = loadQ_io_loadAddrQueue_6; // @[LSQBRAM.scala 144:30:@46680.4]
  assign storeQ_io_loadAddressQueue_7 = loadQ_io_loadAddrQueue_7; // @[LSQBRAM.scala 144:30:@46681.4]
  assign storeQ_io_loadAddressQueue_8 = loadQ_io_loadAddrQueue_8; // @[LSQBRAM.scala 144:30:@46682.4]
  assign storeQ_io_loadAddressQueue_9 = loadQ_io_loadAddrQueue_9; // @[LSQBRAM.scala 144:30:@46683.4]
  assign storeQ_io_loadAddressQueue_10 = loadQ_io_loadAddrQueue_10; // @[LSQBRAM.scala 144:30:@46684.4]
  assign storeQ_io_loadAddressQueue_11 = loadQ_io_loadAddrQueue_11; // @[LSQBRAM.scala 144:30:@46685.4]
  assign storeQ_io_loadAddressQueue_12 = loadQ_io_loadAddrQueue_12; // @[LSQBRAM.scala 144:30:@46686.4]
  assign storeQ_io_loadAddressQueue_13 = loadQ_io_loadAddrQueue_13; // @[LSQBRAM.scala 144:30:@46687.4]
  assign storeQ_io_loadAddressQueue_14 = loadQ_io_loadAddrQueue_14; // @[LSQBRAM.scala 144:30:@46688.4]
  assign storeQ_io_loadAddressQueue_15 = loadQ_io_loadAddrQueue_15; // @[LSQBRAM.scala 144:30:@46689.4]
  assign storeQ_io_storeDataEnable_0 = STORE_DATA_PORT_LSQ_data_io_storeDataEnable; // @[LSQBRAM.scala 156:29:@46791.4]
  assign storeQ_io_dataFromStorePorts_0 = STORE_DATA_PORT_LSQ_data_io_dataToStoreQueue; // @[LSQBRAM.scala 157:32:@46792.4]
  assign storeQ_io_storeAddrEnable_0 = STORE_ADDR_PORT_LSQ_data_io_storeDataEnable; // @[LSQBRAM.scala 158:29:@46793.4]
  assign storeQ_io_addressFromStorePorts_0 = STORE_ADDR_PORT_LSQ_data_io_dataToStoreQueue; // @[LSQBRAM.scala 159:35:@46794.4]
  assign storeQ_io_memIsReadyForStores = io_memIsReadyForStores; // @[LSQBRAM.scala 163:33:@46798.4]
  assign loadQ_clock = clock; // @[:@46335.4]
  assign loadQ_reset = reset; // @[:@46336.4]
  assign loadQ_io_bbStart = GA_io_bbStart; // @[LSQBRAM.scala 113:20:@46540.4]
  assign loadQ_io_bbLoadOffsets_0 = GA_io_bbLoadOffsets_0; // @[LSQBRAM.scala 114:26:@46541.4]
  assign loadQ_io_bbLoadOffsets_1 = GA_io_bbLoadOffsets_1; // @[LSQBRAM.scala 114:26:@46542.4]
  assign loadQ_io_bbLoadOffsets_2 = GA_io_bbLoadOffsets_2; // @[LSQBRAM.scala 114:26:@46543.4]
  assign loadQ_io_bbLoadOffsets_3 = GA_io_bbLoadOffsets_3; // @[LSQBRAM.scala 114:26:@46544.4]
  assign loadQ_io_bbLoadOffsets_4 = GA_io_bbLoadOffsets_4; // @[LSQBRAM.scala 114:26:@46545.4]
  assign loadQ_io_bbLoadOffsets_5 = GA_io_bbLoadOffsets_5; // @[LSQBRAM.scala 114:26:@46546.4]
  assign loadQ_io_bbLoadOffsets_6 = GA_io_bbLoadOffsets_6; // @[LSQBRAM.scala 114:26:@46547.4]
  assign loadQ_io_bbLoadOffsets_7 = GA_io_bbLoadOffsets_7; // @[LSQBRAM.scala 114:26:@46548.4]
  assign loadQ_io_bbLoadOffsets_8 = GA_io_bbLoadOffsets_8; // @[LSQBRAM.scala 114:26:@46549.4]
  assign loadQ_io_bbLoadOffsets_9 = GA_io_bbLoadOffsets_9; // @[LSQBRAM.scala 114:26:@46550.4]
  assign loadQ_io_bbLoadOffsets_10 = GA_io_bbLoadOffsets_10; // @[LSQBRAM.scala 114:26:@46551.4]
  assign loadQ_io_bbLoadOffsets_11 = GA_io_bbLoadOffsets_11; // @[LSQBRAM.scala 114:26:@46552.4]
  assign loadQ_io_bbLoadOffsets_12 = GA_io_bbLoadOffsets_12; // @[LSQBRAM.scala 114:26:@46553.4]
  assign loadQ_io_bbLoadOffsets_13 = GA_io_bbLoadOffsets_13; // @[LSQBRAM.scala 114:26:@46554.4]
  assign loadQ_io_bbLoadOffsets_14 = GA_io_bbLoadOffsets_14; // @[LSQBRAM.scala 114:26:@46555.4]
  assign loadQ_io_bbLoadOffsets_15 = GA_io_bbLoadOffsets_15; // @[LSQBRAM.scala 114:26:@46556.4]
  assign loadQ_io_bbLoadPorts_1 = GA_io_bbLoadPorts_1; // @[LSQBRAM.scala 115:24:@46558.4]
  assign loadQ_io_bbNumLoads = GA_io_bbNumLoads; // @[LSQBRAM.scala 116:23:@46573.4]
  assign loadQ_io_storeTail = storeTail[3:0]; // @[LSQBRAM.scala 106:22:@46473.4]
  assign loadQ_io_storeHead = storeHead[3:0]; // @[LSQBRAM.scala 107:22:@46474.4]
  assign loadQ_io_storeEmpty = storeQ_io_storeEmpty; // @[LSQBRAM.scala 108:23:@46475.4]
  assign loadQ_io_storeAddrDone_0 = storeQ_io_storeAddrDone_0; // @[LSQBRAM.scala 109:26:@46476.4]
  assign loadQ_io_storeAddrDone_1 = storeQ_io_storeAddrDone_1; // @[LSQBRAM.scala 109:26:@46477.4]
  assign loadQ_io_storeAddrDone_2 = storeQ_io_storeAddrDone_2; // @[LSQBRAM.scala 109:26:@46478.4]
  assign loadQ_io_storeAddrDone_3 = storeQ_io_storeAddrDone_3; // @[LSQBRAM.scala 109:26:@46479.4]
  assign loadQ_io_storeAddrDone_4 = storeQ_io_storeAddrDone_4; // @[LSQBRAM.scala 109:26:@46480.4]
  assign loadQ_io_storeAddrDone_5 = storeQ_io_storeAddrDone_5; // @[LSQBRAM.scala 109:26:@46481.4]
  assign loadQ_io_storeAddrDone_6 = storeQ_io_storeAddrDone_6; // @[LSQBRAM.scala 109:26:@46482.4]
  assign loadQ_io_storeAddrDone_7 = storeQ_io_storeAddrDone_7; // @[LSQBRAM.scala 109:26:@46483.4]
  assign loadQ_io_storeAddrDone_8 = storeQ_io_storeAddrDone_8; // @[LSQBRAM.scala 109:26:@46484.4]
  assign loadQ_io_storeAddrDone_9 = storeQ_io_storeAddrDone_9; // @[LSQBRAM.scala 109:26:@46485.4]
  assign loadQ_io_storeAddrDone_10 = storeQ_io_storeAddrDone_10; // @[LSQBRAM.scala 109:26:@46486.4]
  assign loadQ_io_storeAddrDone_11 = storeQ_io_storeAddrDone_11; // @[LSQBRAM.scala 109:26:@46487.4]
  assign loadQ_io_storeAddrDone_12 = storeQ_io_storeAddrDone_12; // @[LSQBRAM.scala 109:26:@46488.4]
  assign loadQ_io_storeAddrDone_13 = storeQ_io_storeAddrDone_13; // @[LSQBRAM.scala 109:26:@46489.4]
  assign loadQ_io_storeAddrDone_14 = storeQ_io_storeAddrDone_14; // @[LSQBRAM.scala 109:26:@46490.4]
  assign loadQ_io_storeAddrDone_15 = storeQ_io_storeAddrDone_15; // @[LSQBRAM.scala 109:26:@46491.4]
  assign loadQ_io_storeDataDone_0 = storeQ_io_storeDataDone_0; // @[LSQBRAM.scala 110:26:@46492.4]
  assign loadQ_io_storeDataDone_1 = storeQ_io_storeDataDone_1; // @[LSQBRAM.scala 110:26:@46493.4]
  assign loadQ_io_storeDataDone_2 = storeQ_io_storeDataDone_2; // @[LSQBRAM.scala 110:26:@46494.4]
  assign loadQ_io_storeDataDone_3 = storeQ_io_storeDataDone_3; // @[LSQBRAM.scala 110:26:@46495.4]
  assign loadQ_io_storeDataDone_4 = storeQ_io_storeDataDone_4; // @[LSQBRAM.scala 110:26:@46496.4]
  assign loadQ_io_storeDataDone_5 = storeQ_io_storeDataDone_5; // @[LSQBRAM.scala 110:26:@46497.4]
  assign loadQ_io_storeDataDone_6 = storeQ_io_storeDataDone_6; // @[LSQBRAM.scala 110:26:@46498.4]
  assign loadQ_io_storeDataDone_7 = storeQ_io_storeDataDone_7; // @[LSQBRAM.scala 110:26:@46499.4]
  assign loadQ_io_storeDataDone_8 = storeQ_io_storeDataDone_8; // @[LSQBRAM.scala 110:26:@46500.4]
  assign loadQ_io_storeDataDone_9 = storeQ_io_storeDataDone_9; // @[LSQBRAM.scala 110:26:@46501.4]
  assign loadQ_io_storeDataDone_10 = storeQ_io_storeDataDone_10; // @[LSQBRAM.scala 110:26:@46502.4]
  assign loadQ_io_storeDataDone_11 = storeQ_io_storeDataDone_11; // @[LSQBRAM.scala 110:26:@46503.4]
  assign loadQ_io_storeDataDone_12 = storeQ_io_storeDataDone_12; // @[LSQBRAM.scala 110:26:@46504.4]
  assign loadQ_io_storeDataDone_13 = storeQ_io_storeDataDone_13; // @[LSQBRAM.scala 110:26:@46505.4]
  assign loadQ_io_storeDataDone_14 = storeQ_io_storeDataDone_14; // @[LSQBRAM.scala 110:26:@46506.4]
  assign loadQ_io_storeDataDone_15 = storeQ_io_storeDataDone_15; // @[LSQBRAM.scala 110:26:@46507.4]
  assign loadQ_io_storeAddrQueue_0 = storeQ_io_storeAddrQueue_0; // @[LSQBRAM.scala 111:27:@46508.4]
  assign loadQ_io_storeAddrQueue_1 = storeQ_io_storeAddrQueue_1; // @[LSQBRAM.scala 111:27:@46509.4]
  assign loadQ_io_storeAddrQueue_2 = storeQ_io_storeAddrQueue_2; // @[LSQBRAM.scala 111:27:@46510.4]
  assign loadQ_io_storeAddrQueue_3 = storeQ_io_storeAddrQueue_3; // @[LSQBRAM.scala 111:27:@46511.4]
  assign loadQ_io_storeAddrQueue_4 = storeQ_io_storeAddrQueue_4; // @[LSQBRAM.scala 111:27:@46512.4]
  assign loadQ_io_storeAddrQueue_5 = storeQ_io_storeAddrQueue_5; // @[LSQBRAM.scala 111:27:@46513.4]
  assign loadQ_io_storeAddrQueue_6 = storeQ_io_storeAddrQueue_6; // @[LSQBRAM.scala 111:27:@46514.4]
  assign loadQ_io_storeAddrQueue_7 = storeQ_io_storeAddrQueue_7; // @[LSQBRAM.scala 111:27:@46515.4]
  assign loadQ_io_storeAddrQueue_8 = storeQ_io_storeAddrQueue_8; // @[LSQBRAM.scala 111:27:@46516.4]
  assign loadQ_io_storeAddrQueue_9 = storeQ_io_storeAddrQueue_9; // @[LSQBRAM.scala 111:27:@46517.4]
  assign loadQ_io_storeAddrQueue_10 = storeQ_io_storeAddrQueue_10; // @[LSQBRAM.scala 111:27:@46518.4]
  assign loadQ_io_storeAddrQueue_11 = storeQ_io_storeAddrQueue_11; // @[LSQBRAM.scala 111:27:@46519.4]
  assign loadQ_io_storeAddrQueue_12 = storeQ_io_storeAddrQueue_12; // @[LSQBRAM.scala 111:27:@46520.4]
  assign loadQ_io_storeAddrQueue_13 = storeQ_io_storeAddrQueue_13; // @[LSQBRAM.scala 111:27:@46521.4]
  assign loadQ_io_storeAddrQueue_14 = storeQ_io_storeAddrQueue_14; // @[LSQBRAM.scala 111:27:@46522.4]
  assign loadQ_io_storeAddrQueue_15 = storeQ_io_storeAddrQueue_15; // @[LSQBRAM.scala 111:27:@46523.4]
  assign loadQ_io_storeDataQueue_0 = storeQ_io_storeDataQueue_0; // @[LSQBRAM.scala 112:27:@46524.4]
  assign loadQ_io_storeDataQueue_1 = storeQ_io_storeDataQueue_1; // @[LSQBRAM.scala 112:27:@46525.4]
  assign loadQ_io_storeDataQueue_2 = storeQ_io_storeDataQueue_2; // @[LSQBRAM.scala 112:27:@46526.4]
  assign loadQ_io_storeDataQueue_3 = storeQ_io_storeDataQueue_3; // @[LSQBRAM.scala 112:27:@46527.4]
  assign loadQ_io_storeDataQueue_4 = storeQ_io_storeDataQueue_4; // @[LSQBRAM.scala 112:27:@46528.4]
  assign loadQ_io_storeDataQueue_5 = storeQ_io_storeDataQueue_5; // @[LSQBRAM.scala 112:27:@46529.4]
  assign loadQ_io_storeDataQueue_6 = storeQ_io_storeDataQueue_6; // @[LSQBRAM.scala 112:27:@46530.4]
  assign loadQ_io_storeDataQueue_7 = storeQ_io_storeDataQueue_7; // @[LSQBRAM.scala 112:27:@46531.4]
  assign loadQ_io_storeDataQueue_8 = storeQ_io_storeDataQueue_8; // @[LSQBRAM.scala 112:27:@46532.4]
  assign loadQ_io_storeDataQueue_9 = storeQ_io_storeDataQueue_9; // @[LSQBRAM.scala 112:27:@46533.4]
  assign loadQ_io_storeDataQueue_10 = storeQ_io_storeDataQueue_10; // @[LSQBRAM.scala 112:27:@46534.4]
  assign loadQ_io_storeDataQueue_11 = storeQ_io_storeDataQueue_11; // @[LSQBRAM.scala 112:27:@46535.4]
  assign loadQ_io_storeDataQueue_12 = storeQ_io_storeDataQueue_12; // @[LSQBRAM.scala 112:27:@46536.4]
  assign loadQ_io_storeDataQueue_13 = storeQ_io_storeDataQueue_13; // @[LSQBRAM.scala 112:27:@46537.4]
  assign loadQ_io_storeDataQueue_14 = storeQ_io_storeDataQueue_14; // @[LSQBRAM.scala 112:27:@46538.4]
  assign loadQ_io_storeDataQueue_15 = storeQ_io_storeDataQueue_15; // @[LSQBRAM.scala 112:27:@46539.4]
  assign loadQ_io_loadAddrEnable_0 = LOAD_PORT_LSQ_data_io_loadAddrEnable; // @[LSQBRAM.scala 130:32:@46629.4]
  assign loadQ_io_loadAddrEnable_1 = LOAD_PORT_LSQ_data_1_io_loadAddrEnable; // @[LSQBRAM.scala 130:32:@46634.4]
  assign loadQ_io_addrFromLoadPorts_0 = LOAD_PORT_LSQ_data_io_addrToLoadQueue; // @[LSQBRAM.scala 129:35:@46628.4]
  assign loadQ_io_addrFromLoadPorts_1 = LOAD_PORT_LSQ_data_1_io_addrToLoadQueue; // @[LSQBRAM.scala 129:35:@46633.4]
  assign loadQ_io_loadPorts_0_ready = LOAD_PORT_LSQ_data_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 127:33:@46627.4]
  assign loadQ_io_loadPorts_1_ready = LOAD_PORT_LSQ_data_1_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 127:33:@46632.4]
  assign loadQ_io_loadDataFromMem = io_loadDataIn; // @[LSQBRAM.scala 133:28:@46635.4]
  assign loadQ_io_memIsReadyForLoads = io_memIsReadyForLoads; // @[LSQBRAM.scala 134:31:@46636.4]
  assign GA_io_loadTail = loadTail[3:0]; // @[LSQBRAM.scala 91:18:@46426.4]
  assign GA_io_loadHead = loadHead[3:0]; // @[LSQBRAM.scala 92:18:@46427.4]
  assign GA_io_loadEmpty = loadQ_io_loadEmpty; // @[LSQBRAM.scala 93:19:@46428.4]
  assign GA_io_storeTail = storeTail[3:0]; // @[LSQBRAM.scala 97:19:@46462.4]
  assign GA_io_storeHead = storeHead[3:0]; // @[LSQBRAM.scala 98:19:@46463.4]
  assign GA_io_storeEmpty = storeQ_io_storeEmpty; // @[LSQBRAM.scala 99:20:@46464.4]
  assign GA_io_bbStartSignals_0 = io_bbpValids_0; // @[LSQBRAM.scala 101:24:@46466.4]
  assign GA_io_bbStartSignals_1 = io_bbpValids_1; // @[LSQBRAM.scala 101:24:@46467.4]
  assign LOAD_PORT_LSQ_data_clock = clock; // @[:@46341.4]
  assign LOAD_PORT_LSQ_data_reset = reset; // @[:@46342.4]
  assign LOAD_PORT_LSQ_data_io_addrFromPrev_valid = io_rdPortsPrev_0_valid; // @[LSQBRAM.scala 76:26:@46357.4]
  assign LOAD_PORT_LSQ_data_io_addrFromPrev_bits = io_rdPortsPrev_0_bits; // @[LSQBRAM.scala 76:26:@46356.4]
  assign LOAD_PORT_LSQ_data_io_portEnable = GA_io_loadPortsEnable_0; // @[LSQBRAM.scala 76:26:@46355.4]
  assign LOAD_PORT_LSQ_data_io_dataToNext_ready = io_rdPortsNext_0_ready; // @[LSQBRAM.scala 76:26:@46354.4]
  assign LOAD_PORT_LSQ_data_io_dataFromLoadQueue_valid = loadQ_io_loadPorts_0_valid; // @[LSQBRAM.scala 76:26:@46348.4]
  assign LOAD_PORT_LSQ_data_io_dataFromLoadQueue_bits = loadQ_io_loadPorts_0_bits; // @[LSQBRAM.scala 76:26:@46347.4]
  assign LOAD_PORT_LSQ_data_1_clock = clock; // @[:@46344.4]
  assign LOAD_PORT_LSQ_data_1_reset = reset; // @[:@46345.4]
  assign LOAD_PORT_LSQ_data_1_io_addrFromPrev_valid = io_rdPortsPrev_1_valid; // @[LSQBRAM.scala 76:26:@46369.4]
  assign LOAD_PORT_LSQ_data_1_io_addrFromPrev_bits = io_rdPortsPrev_1_bits; // @[LSQBRAM.scala 76:26:@46368.4]
  assign LOAD_PORT_LSQ_data_1_io_portEnable = GA_io_loadPortsEnable_1; // @[LSQBRAM.scala 76:26:@46367.4]
  assign LOAD_PORT_LSQ_data_1_io_dataToNext_ready = io_rdPortsNext_1_ready; // @[LSQBRAM.scala 76:26:@46366.4]
  assign LOAD_PORT_LSQ_data_1_io_dataFromLoadQueue_valid = loadQ_io_loadPorts_1_valid; // @[LSQBRAM.scala 76:26:@46360.4]
  assign LOAD_PORT_LSQ_data_1_io_dataFromLoadQueue_bits = loadQ_io_loadPorts_1_bits; // @[LSQBRAM.scala 76:26:@46359.4]
  assign STORE_DATA_PORT_LSQ_data_clock = clock; // @[:@46372.4]
  assign STORE_DATA_PORT_LSQ_data_reset = reset; // @[:@46373.4]
  assign STORE_DATA_PORT_LSQ_data_io_dataFromPrev_valid = io_wrDataPorts_0_valid; // @[LSQBRAM.scala 79:31:@46379.4]
  assign STORE_DATA_PORT_LSQ_data_io_dataFromPrev_bits = io_wrDataPorts_0_bits; // @[LSQBRAM.scala 79:31:@46378.4]
  assign STORE_DATA_PORT_LSQ_data_io_portEnable = GA_io_storePortsEnable_0; // @[LSQBRAM.scala 79:31:@46377.4]
  assign STORE_ADDR_PORT_LSQ_data_clock = clock; // @[:@46382.4]
  assign STORE_ADDR_PORT_LSQ_data_reset = reset; // @[:@46383.4]
  assign STORE_ADDR_PORT_LSQ_data_io_dataFromPrev_valid = io_wrAddrPorts_0_valid; // @[LSQBRAM.scala 82:34:@46389.4]
  assign STORE_ADDR_PORT_LSQ_data_io_dataFromPrev_bits = io_wrAddrPorts_0_bits; // @[LSQBRAM.scala 82:34:@46388.4]
  assign STORE_ADDR_PORT_LSQ_data_io_portEnable = GA_io_storePortsEnable_0; // @[LSQBRAM.scala 82:34:@46387.4]
endmodule
